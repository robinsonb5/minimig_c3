-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity DiagROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end DiagROM_ROM;

architecture arch of DiagROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ed040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"880d8004",
     5 => x"84808080",
     6 => x"940471fd",
     7 => x"06087283",
     8 => x"06098105",
     9 => x"8205832b",
    10 => x"2a83ffff",
    11 => x"06520471",
    12 => x"fc060872",
    13 => x"83060981",
    14 => x"05830510",
    15 => x"10102a81",
    16 => x"ff065204",
    17 => x"71fc0608",
    18 => x"8480809f",
    19 => x"d8738306",
    20 => x"10100508",
    21 => x"067381ff",
    22 => x"06738306",
    23 => x"09810583",
    24 => x"05101010",
    25 => x"2b0772fc",
    26 => x"060c5151",
    27 => x"04028405",
    28 => x"84808080",
    29 => x"880c8480",
    30 => x"8080940b",
    31 => x"8480808f",
    32 => x"da040000",
    33 => x"02c4050d",
    34 => x"0280c005",
    35 => x"9fe0e05b",
    36 => x"56807670",
    37 => x"84055808",
    38 => x"715e5e57",
    39 => x"7c708405",
    40 => x"5e085880",
    41 => x"5b77982a",
    42 => x"78882b59",
    43 => x"54738938",
    44 => x"765e8480",
    45 => x"8083e204",
    46 => x"7b802e81",
    47 => x"fd38805c",
    48 => x"7380e42e",
    49 => x"a1387380",
    50 => x"e4268e38",
    51 => x"7380e32e",
    52 => x"819a3884",
    53 => x"808082fa",
    54 => x"047380f3",
    55 => x"2e80f538",
    56 => x"84808082",
    57 => x"fa047584",
    58 => x"1771087e",
    59 => x"5c555752",
    60 => x"7280258e",
    61 => x"38ad5184",
    62 => x"80808fcc",
    63 => x"2d720981",
    64 => x"05537280",
    65 => x"2ebe3887",
    66 => x"55729c2a",
    67 => x"73842b54",
    68 => x"5271802e",
    69 => x"83388159",
    70 => x"8972258a",
    71 => x"38b71252",
    72 => x"84808082",
    73 => x"a904b012",
    74 => x"5278802e",
    75 => x"89387151",
    76 => x"8480808f",
    77 => x"cc2dff15",
    78 => x"55748025",
    79 => x"cc388480",
    80 => x"8082cc04",
    81 => x"b0518480",
    82 => x"808fcc2d",
    83 => x"80538480",
    84 => x"80839304",
    85 => x"75841771",
    86 => x"0870545c",
    87 => x"57528480",
    88 => x"8085ab2d",
    89 => x"7b538480",
    90 => x"80839304",
    91 => x"75841771",
    92 => x"08565752",
    93 => x"84808083",
    94 => x"ca04a551",
    95 => x"8480808f",
    96 => x"cc2d7351",
    97 => x"8480808f",
    98 => x"cc2d8217",
    99 => x"57848080",
   100 => x"83d50472",
   101 => x"ff145452",
   102 => x"807225b9",
   103 => x"38797081",
   104 => x"055b8480",
   105 => x"8080af2d",
   106 => x"70525484",
   107 => x"80808fcc",
   108 => x"2d811757",
   109 => x"84808083",
   110 => x"930473a5",
   111 => x"2e098106",
   112 => x"8938815c",
   113 => x"84808083",
   114 => x"d5047351",
   115 => x"8480808f",
   116 => x"cc2d8117",
   117 => x"57811b5b",
   118 => x"837b25fd",
   119 => x"c83873fd",
   120 => x"bb387d9f",
   121 => x"e0800c02",
   122 => x"bc050d04",
   123 => x"02f4050d",
   124 => x"7470882a",
   125 => x"83fe8006",
   126 => x"7072982a",
   127 => x"0772882b",
   128 => x"87fc8080",
   129 => x"0673982b",
   130 => x"81f00a06",
   131 => x"71730707",
   132 => x"9fe0800c",
   133 => x"56515351",
   134 => x"028c050d",
   135 => x"0402f805",
   136 => x"0d028e05",
   137 => x"84808080",
   138 => x"af2d7498",
   139 => x"2b71902b",
   140 => x"0770902c",
   141 => x"9fe0800c",
   142 => x"52520288",
   143 => x"050d0402",
   144 => x"f8050d73",
   145 => x"70902b71",
   146 => x"902a079f",
   147 => x"e0800c52",
   148 => x"0288050d",
   149 => x"0402f805",
   150 => x"0d735170",
   151 => x"802e8c38",
   152 => x"709fe1a0",
   153 => x"0c800b9f",
   154 => x"e1a80c9f",
   155 => x"e1a80852",
   156 => x"7198389f",
   157 => x"e1a00884",
   158 => x"119fe1a0",
   159 => x"0c70089f",
   160 => x"e1a40c51",
   161 => x"84808085",
   162 => x"94049fe1",
   163 => x"a408882b",
   164 => x"9fe1a40c",
   165 => x"81128306",
   166 => x"9fe1a80c",
   167 => x"9fe1a408",
   168 => x"982c9fe0",
   169 => x"800c0288",
   170 => x"050d0402",
   171 => x"e8050d77",
   172 => x"70525684",
   173 => x"808084d5",
   174 => x"2d9fe080",
   175 => x"08528053",
   176 => x"71802e97",
   177 => x"38811353",
   178 => x"80518480",
   179 => x"8084d52d",
   180 => x"9fe08008",
   181 => x"52848080",
   182 => x"85c00482",
   183 => x"13548155",
   184 => x"900b86e9",
   185 => x"808423a0",
   186 => x"810b86e9",
   187 => x"80802386",
   188 => x"e9808022",
   189 => x"52800b86",
   190 => x"e9808023",
   191 => x"86e98080",
   192 => x"2253800b",
   193 => x"86e98080",
   194 => x"2386e980",
   195 => x"80227083",
   196 => x"ffff0673",
   197 => x"882a7081",
   198 => x"06515451",
   199 => x"5371802e",
   200 => x"81a43874",
   201 => x"802e80e0",
   202 => x"38728280",
   203 => x"862e0981",
   204 => x"06819338",
   205 => x"8055fed5",
   206 => x"ca0b86e9",
   207 => x"80802386",
   208 => x"e9808022",
   209 => x"52810b86",
   210 => x"e9808023",
   211 => x"86e98080",
   212 => x"22527486",
   213 => x"e9808023",
   214 => x"86e98080",
   215 => x"22527386",
   216 => x"e9808023",
   217 => x"86e98080",
   218 => x"22527486",
   219 => x"e9808023",
   220 => x"86e98080",
   221 => x"22527486",
   222 => x"e9808023",
   223 => x"86e98080",
   224 => x"22528480",
   225 => x"8087c604",
   226 => x"73812a82",
   227 => x"80800752",
   228 => x"72722e09",
   229 => x"8106af38",
   230 => x"75518480",
   231 => x"8084d52d",
   232 => x"9fe08008",
   233 => x"53ff1454",
   234 => x"73ff2ea7",
   235 => x"387286e9",
   236 => x"80803486",
   237 => x"e9808033",
   238 => x"5272802e",
   239 => x"e8388051",
   240 => x"84808087",
   241 => x"9a04910b",
   242 => x"86e98084",
   243 => x"23848080",
   244 => x"85e00491",
   245 => x"0b86e980",
   246 => x"8423810b",
   247 => x"9fe0800c",
   248 => x"0298050d",
   249 => x"0402f405",
   250 => x"0d86e980",
   251 => x"805281ff",
   252 => x"72237122",
   253 => x"5381ff72",
   254 => x"2372882b",
   255 => x"83fe8006",
   256 => x"72227081",
   257 => x"ff065152",
   258 => x"5381ff72",
   259 => x"23727107",
   260 => x"882b7222",
   261 => x"7081ff06",
   262 => x"51525381",
   263 => x"ff722372",
   264 => x"7107882b",
   265 => x"72227081",
   266 => x"ff067207",
   267 => x"9fe0800c",
   268 => x"5253028c",
   269 => x"050d0402",
   270 => x"f4050d74",
   271 => x"767181ff",
   272 => x"06535353",
   273 => x"7086e980",
   274 => x"80239fe1",
   275 => x"ac088538",
   276 => x"71892b52",
   277 => x"71982a51",
   278 => x"7086e980",
   279 => x"80237190",
   280 => x"2a7081ff",
   281 => x"06515170",
   282 => x"86e98080",
   283 => x"2371882a",
   284 => x"7081ff06",
   285 => x"51517086",
   286 => x"e9808023",
   287 => x"7181ff06",
   288 => x"517086e9",
   289 => x"80802372",
   290 => x"902a7081",
   291 => x"ff065151",
   292 => x"7086e980",
   293 => x"802386e9",
   294 => x"80802270",
   295 => x"81ff0651",
   296 => x"5182b8bf",
   297 => x"527081ff",
   298 => x"2e098106",
   299 => x"9a3881ff",
   300 => x"0b86e980",
   301 => x"802386e9",
   302 => x"80802270",
   303 => x"81ff06ff",
   304 => x"14545151",
   305 => x"71df3870",
   306 => x"9fe0800c",
   307 => x"028c050d",
   308 => x"0402fc05",
   309 => x"0d81c751",
   310 => x"81ff0b86",
   311 => x"e9808023",
   312 => x"ff115170",
   313 => x"8025f138",
   314 => x"0284050d",
   315 => x"0402f005",
   316 => x"0d848080",
   317 => x"89d12d81",
   318 => x"9c9f5380",
   319 => x"5287fc80",
   320 => x"f7518480",
   321 => x"8088b72d",
   322 => x"9fe08008",
   323 => x"549fe080",
   324 => x"08812e09",
   325 => x"8106b338",
   326 => x"81ff0b86",
   327 => x"e9808023",
   328 => x"820a5284",
   329 => x"9c80e951",
   330 => x"84808088",
   331 => x"b72d9fe0",
   332 => x"80089138",
   333 => x"81ff0b86",
   334 => x"e9808023",
   335 => x"73538480",
   336 => x"808ad104",
   337 => x"84808089",
   338 => x"d12dff13",
   339 => x"5372ffab",
   340 => x"38729fe0",
   341 => x"800c0290",
   342 => x"050d0402",
   343 => x"f4050d81",
   344 => x"ff0b86e9",
   345 => x"80802384",
   346 => x"80809fe8",
   347 => x"51848080",
   348 => x"85ab2d93",
   349 => x"53805287",
   350 => x"fc80c151",
   351 => x"84808088",
   352 => x"b72d9fe0",
   353 => x"80089138",
   354 => x"81ff0b86",
   355 => x"e9808023",
   356 => x"81538480",
   357 => x"808ba404",
   358 => x"84808089",
   359 => x"d12dff13",
   360 => x"5372d238",
   361 => x"729fe080",
   362 => x"0c028c05",
   363 => x"0d0402f0",
   364 => x"050d8480",
   365 => x"8089d12d",
   366 => x"83aa5284",
   367 => x"9c80c851",
   368 => x"84808088",
   369 => x"b72d9fe0",
   370 => x"8008812e",
   371 => x"09810696",
   372 => x"38848080",
   373 => x"87e52d9f",
   374 => x"e0800883",
   375 => x"ffff0653",
   376 => x"7283aa2e",
   377 => x"9d388480",
   378 => x"808adb2d",
   379 => x"8480808b",
   380 => x"fa048154",
   381 => x"8480808d",
   382 => x"84048054",
   383 => x"8480808d",
   384 => x"840481ff",
   385 => x"0b86e980",
   386 => x"8023b153",
   387 => x"84808089",
   388 => x"ed2d9fe0",
   389 => x"8008802e",
   390 => x"80db3880",
   391 => x"5287fc80",
   392 => x"fa518480",
   393 => x"8088b72d",
   394 => x"9fe08008",
   395 => x"80c73881",
   396 => x"ff0b86e9",
   397 => x"80802386",
   398 => x"e9808022",
   399 => x"5381ff0b",
   400 => x"86e98080",
   401 => x"2381ff0b",
   402 => x"86e98080",
   403 => x"2381ff0b",
   404 => x"86e98080",
   405 => x"2381ff0b",
   406 => x"86e98080",
   407 => x"2372862a",
   408 => x"7081069f",
   409 => x"e0800856",
   410 => x"51537280",
   411 => x"2e963884",
   412 => x"80808bf2",
   413 => x"0472822e",
   414 => x"ff8038ff",
   415 => x"135372ff",
   416 => x"8b387254",
   417 => x"739fe080",
   418 => x"0c029005",
   419 => x"0d0402f4",
   420 => x"050d810b",
   421 => x"9fe1ac0c",
   422 => x"a00b86e9",
   423 => x"80882383",
   424 => x"0b86e980",
   425 => x"84238480",
   426 => x"8089d12d",
   427 => x"820b86e9",
   428 => x"80842387",
   429 => x"53805284",
   430 => x"d480c051",
   431 => x"84808088",
   432 => x"b72d9fe0",
   433 => x"8008812e",
   434 => x"97387282",
   435 => x"2e098106",
   436 => x"89388053",
   437 => x"8480808e",
   438 => x"9404ff13",
   439 => x"5372d638",
   440 => x"8480808b",
   441 => x"ae2d9fe0",
   442 => x"80089fe1",
   443 => x"ac0c8152",
   444 => x"87fc80d0",
   445 => x"51848080",
   446 => x"88b72d81",
   447 => x"ff0b86e9",
   448 => x"80802383",
   449 => x"0b86e980",
   450 => x"842381ff",
   451 => x"0b86e980",
   452 => x"80238153",
   453 => x"729fe080",
   454 => x"0c028c05",
   455 => x"0d04800b",
   456 => x"9fe0800c",
   457 => x"0402e805",
   458 => x"0d785680",
   459 => x"5581ff0b",
   460 => x"86e98080",
   461 => x"23820b86",
   462 => x"e9808423",
   463 => x"810b86e9",
   464 => x"80882381",
   465 => x"ff0b86e9",
   466 => x"80802377",
   467 => x"5287fc80",
   468 => x"d1518480",
   469 => x"8088b72d",
   470 => x"74539fe0",
   471 => x"8008752e",
   472 => x"09810680",
   473 => x"dd3880db",
   474 => x"c6df5481",
   475 => x"ff0b86e9",
   476 => x"80802386",
   477 => x"e9808022",
   478 => x"7081ff06",
   479 => x"51537281",
   480 => x"fe2e0981",
   481 => x"06a43880",
   482 => x"ff538480",
   483 => x"8087e52d",
   484 => x"9fe08008",
   485 => x"76708405",
   486 => x"580cff13",
   487 => x"53728025",
   488 => x"e9388155",
   489 => x"8480808f",
   490 => x"b104ff14",
   491 => x"5473ffbb",
   492 => x"3881ff0b",
   493 => x"86e98080",
   494 => x"23830b86",
   495 => x"e9808423",
   496 => x"7453729f",
   497 => x"e0800c02",
   498 => x"98050d04",
   499 => x"02fc050d",
   500 => x"709fe080",
   501 => x"0c028405",
   502 => x"0d0402f8",
   503 => x"050d8480",
   504 => x"809ff451",
   505 => x"84808085",
   506 => x"ab2d8480",
   507 => x"808d8e2d",
   508 => x"9fe08008",
   509 => x"802ebb38",
   510 => x"848080a0",
   511 => x"8c518480",
   512 => x"8085ab2d",
   513 => x"84808091",
   514 => x"942d8052",
   515 => x"848080a0",
   516 => x"a4518480",
   517 => x"809d8b2d",
   518 => x"9fe08008",
   519 => x"802e8738",
   520 => x"84808080",
   521 => x"8c2d8480",
   522 => x"80a0b051",
   523 => x"84808085",
   524 => x"ab2d8480",
   525 => x"80a0c851",
   526 => x"84808085",
   527 => x"ab2d800b",
   528 => x"9fe0800c",
   529 => x"0288050d",
   530 => x"0402e805",
   531 => x"0d77797b",
   532 => x"58555580",
   533 => x"53727625",
   534 => x"af387470",
   535 => x"81055684",
   536 => x"808080af",
   537 => x"2d747081",
   538 => x"05568480",
   539 => x"8080af2d",
   540 => x"52527171",
   541 => x"2e893881",
   542 => x"51848080",
   543 => x"918a0481",
   544 => x"13538480",
   545 => x"8090d504",
   546 => x"8051709f",
   547 => x"e0800c02",
   548 => x"98050d04",
   549 => x"02d8050d",
   550 => x"ff0b9fe5",
   551 => x"d80c800b",
   552 => x"9fe5ec0c",
   553 => x"848080a0",
   554 => x"e8518480",
   555 => x"8085ab2d",
   556 => x"9fe1c452",
   557 => x"80518480",
   558 => x"808ea52d",
   559 => x"9fe08008",
   560 => x"549fe080",
   561 => x"08953884",
   562 => x"8080a0f8",
   563 => x"51848080",
   564 => x"85ab2d73",
   565 => x"55848080",
   566 => x"98ef0484",
   567 => x"8080a18c",
   568 => x"51848080",
   569 => x"85ab2d80",
   570 => x"56810b9f",
   571 => x"e1b80c88",
   572 => x"53848080",
   573 => x"a1a4529f",
   574 => x"e1fa5184",
   575 => x"808090c9",
   576 => x"2d9fe080",
   577 => x"08762e09",
   578 => x"81068938",
   579 => x"9fe08008",
   580 => x"9fe1b80c",
   581 => x"88538480",
   582 => x"80a1b052",
   583 => x"9fe29651",
   584 => x"84808090",
   585 => x"c92d9fe0",
   586 => x"80088938",
   587 => x"9fe08008",
   588 => x"9fe1b80c",
   589 => x"9fe1b808",
   590 => x"52848080",
   591 => x"a1bc5184",
   592 => x"80808184",
   593 => x"2d9fe1b8",
   594 => x"08802e81",
   595 => x"c1389fe5",
   596 => x"8a0b8480",
   597 => x"8080af2d",
   598 => x"9fe58b0b",
   599 => x"84808080",
   600 => x"af2d7198",
   601 => x"2b71902b",
   602 => x"079fe58c",
   603 => x"0b848080",
   604 => x"80af2d70",
   605 => x"882b7207",
   606 => x"9fe58d0b",
   607 => x"84808080",
   608 => x"af2d7107",
   609 => x"9fe5c20b",
   610 => x"84808080",
   611 => x"af2d9fe5",
   612 => x"c30b8480",
   613 => x"8080af2d",
   614 => x"71882b07",
   615 => x"535f5452",
   616 => x"5a565755",
   617 => x"7381abaa",
   618 => x"2e098106",
   619 => x"94387551",
   620 => x"84808083",
   621 => x"ec2d9fe0",
   622 => x"80085684",
   623 => x"808093da",
   624 => x"047382d4",
   625 => x"d52e9338",
   626 => x"848080a1",
   627 => x"d0518480",
   628 => x"8085ab2d",
   629 => x"84808095",
   630 => x"d9047552",
   631 => x"848080a1",
   632 => x"f0518480",
   633 => x"8081842d",
   634 => x"9fe1c452",
   635 => x"75518480",
   636 => x"808ea52d",
   637 => x"9fe08008",
   638 => x"559fe080",
   639 => x"08802e84",
   640 => x"ee388480",
   641 => x"80a28851",
   642 => x"84808085",
   643 => x"ab2d8480",
   644 => x"80a2b051",
   645 => x"84808081",
   646 => x"842d8853",
   647 => x"848080a1",
   648 => x"b0529fe2",
   649 => x"96518480",
   650 => x"8090c92d",
   651 => x"9fe08008",
   652 => x"8d38810b",
   653 => x"9fe5ec0c",
   654 => x"84808094",
   655 => x"ea048853",
   656 => x"848080a1",
   657 => x"a4529fe1",
   658 => x"fa518480",
   659 => x"8090c92d",
   660 => x"9fe08008",
   661 => x"802e9338",
   662 => x"848080a2",
   663 => x"c8518480",
   664 => x"8081842d",
   665 => x"84808095",
   666 => x"d9049fe5",
   667 => x"c20b8480",
   668 => x"8080af2d",
   669 => x"547380d5",
   670 => x"2e098106",
   671 => x"80db389f",
   672 => x"e5c30b84",
   673 => x"808080af",
   674 => x"2d547381",
   675 => x"aa2e0981",
   676 => x"0680c638",
   677 => x"800b9fe1",
   678 => x"c40b8480",
   679 => x"8080af2d",
   680 => x"56547481",
   681 => x"e92e8338",
   682 => x"81547481",
   683 => x"eb2e8c38",
   684 => x"80557375",
   685 => x"2e098106",
   686 => x"83b5389f",
   687 => x"e1cf0b84",
   688 => x"808080af",
   689 => x"2d557491",
   690 => x"389fe1d0",
   691 => x"0b848080",
   692 => x"80af2d54",
   693 => x"73822e89",
   694 => x"38805584",
   695 => x"808098ef",
   696 => x"049fe1d1",
   697 => x"0b848080",
   698 => x"80af2d70",
   699 => x"9fe5f40c",
   700 => x"ff059fe5",
   701 => x"e80c9fe1",
   702 => x"d20b8480",
   703 => x"8080af2d",
   704 => x"9fe1d30b",
   705 => x"84808080",
   706 => x"af2d5876",
   707 => x"05778280",
   708 => x"2905709f",
   709 => x"e5dc0c9f",
   710 => x"e1d40b84",
   711 => x"808080af",
   712 => x"2d709fe5",
   713 => x"d40c9fe5",
   714 => x"ec085957",
   715 => x"5876802e",
   716 => x"81d73888",
   717 => x"53848080",
   718 => x"a1b0529f",
   719 => x"e2965184",
   720 => x"808090c9",
   721 => x"2d9fe080",
   722 => x"0882a438",
   723 => x"9fe5f408",
   724 => x"70842b9f",
   725 => x"e5c40c70",
   726 => x"9fe5f00c",
   727 => x"9fe1e90b",
   728 => x"84808080",
   729 => x"af2d9fe1",
   730 => x"e80b8480",
   731 => x"8080af2d",
   732 => x"71828029",
   733 => x"059fe1ea",
   734 => x"0b848080",
   735 => x"80af2d70",
   736 => x"84808029",
   737 => x"129fe1eb",
   738 => x"0b848080",
   739 => x"80af2d70",
   740 => x"81800a29",
   741 => x"12709fe1",
   742 => x"bc0c9fe5",
   743 => x"d4087129",
   744 => x"9fe5dc08",
   745 => x"05709fe5",
   746 => x"fc0c9fe1",
   747 => x"f10b8480",
   748 => x"8080af2d",
   749 => x"9fe1f00b",
   750 => x"84808080",
   751 => x"af2d7182",
   752 => x"8029059f",
   753 => x"e1f20b84",
   754 => x"808080af",
   755 => x"2d708480",
   756 => x"8029129f",
   757 => x"e1f30b84",
   758 => x"808080af",
   759 => x"2d70982b",
   760 => x"81f00a06",
   761 => x"7205709f",
   762 => x"e1c00cfe",
   763 => x"117e2977",
   764 => x"059fe5e4",
   765 => x"0c525952",
   766 => x"43545e51",
   767 => x"5259525d",
   768 => x"57595784",
   769 => x"808098ed",
   770 => x"049fe1d6",
   771 => x"0b848080",
   772 => x"80af2d9f",
   773 => x"e1d50b84",
   774 => x"808080af",
   775 => x"2d718280",
   776 => x"2905709f",
   777 => x"e5c40c70",
   778 => x"a02983ff",
   779 => x"0570892a",
   780 => x"709fe5f0",
   781 => x"0c9fe1db",
   782 => x"0b848080",
   783 => x"80af2d9f",
   784 => x"e1da0b84",
   785 => x"808080af",
   786 => x"2d718280",
   787 => x"2905709f",
   788 => x"e1bc0c7b",
   789 => x"71291e70",
   790 => x"9fe5e40c",
   791 => x"7d9fe1c0",
   792 => x"0c73059f",
   793 => x"e5fc0c55",
   794 => x"5e515155",
   795 => x"55815574",
   796 => x"9fe0800c",
   797 => x"02a8050d",
   798 => x"0402ec05",
   799 => x"0d767087",
   800 => x"2c7180ff",
   801 => x"06575553",
   802 => x"9fe5ec08",
   803 => x"8a387288",
   804 => x"2c7381ff",
   805 => x"06565473",
   806 => x"9fe5d808",
   807 => x"2ea4389f",
   808 => x"e1c4529f",
   809 => x"e5dc0814",
   810 => x"51848080",
   811 => x"8ea52d9f",
   812 => x"e0800853",
   813 => x"9fe08008",
   814 => x"802e80c9",
   815 => x"38739fe5",
   816 => x"d80c9fe5",
   817 => x"ec08802e",
   818 => x"a0387484",
   819 => x"299fe1c4",
   820 => x"05700852",
   821 => x"53848080",
   822 => x"83ec2d9f",
   823 => x"e08008f0",
   824 => x"0a065584",
   825 => x"80809a83",
   826 => x"0474109f",
   827 => x"e1c40570",
   828 => x"84808080",
   829 => x"9a2d5253",
   830 => x"84808084",
   831 => x"9d2d9fe0",
   832 => x"80085574",
   833 => x"53729fe0",
   834 => x"800c0294",
   835 => x"050d0402",
   836 => x"cc050d7e",
   837 => x"605e5b80",
   838 => x"56ff0b9f",
   839 => x"e5d80c9f",
   840 => x"e1c0089f",
   841 => x"e5e40856",
   842 => x"579fe5ec",
   843 => x"08762e8e",
   844 => x"389fe5f4",
   845 => x"08842b59",
   846 => x"8480809a",
   847 => x"c5049fe5",
   848 => x"f008842b",
   849 => x"59805a79",
   850 => x"792781e8",
   851 => x"38798f06",
   852 => x"a0175754",
   853 => x"73a23874",
   854 => x"52848080",
   855 => x"a2e85184",
   856 => x"80808184",
   857 => x"2d9fe1c4",
   858 => x"52745181",
   859 => x"15558480",
   860 => x"808ea52d",
   861 => x"9fe1c456",
   862 => x"80768480",
   863 => x"8080af2d",
   864 => x"55587378",
   865 => x"2e833881",
   866 => x"587381e5",
   867 => x"2e819c38",
   868 => x"81707906",
   869 => x"555c7380",
   870 => x"2e819038",
   871 => x"8b168480",
   872 => x"8080af2d",
   873 => x"98065877",
   874 => x"8181388b",
   875 => x"537c5275",
   876 => x"51848080",
   877 => x"90c92d9f",
   878 => x"e0800880",
   879 => x"ee389c16",
   880 => x"08518480",
   881 => x"8083ec2d",
   882 => x"9fe08008",
   883 => x"841c0c9a",
   884 => x"16848080",
   885 => x"809a2d51",
   886 => x"84808084",
   887 => x"9d2d9fe0",
   888 => x"80089fe0",
   889 => x"80085555",
   890 => x"9fe5ec08",
   891 => x"802e9f38",
   892 => x"94168480",
   893 => x"80809a2d",
   894 => x"51848080",
   895 => x"849d2d9f",
   896 => x"e0800890",
   897 => x"2b83fff0",
   898 => x"0a067016",
   899 => x"51547388",
   900 => x"1c0c777b",
   901 => x"0c7c5284",
   902 => x"8080a388",
   903 => x"51848080",
   904 => x"81842d7b",
   905 => x"54848080",
   906 => x"9d810481",
   907 => x"1a5a8480",
   908 => x"809ac704",
   909 => x"9fe5ec08",
   910 => x"802e80c3",
   911 => x"38765184",
   912 => x"808098f9",
   913 => x"2d9fe080",
   914 => x"089fe080",
   915 => x"08538480",
   916 => x"80a39c52",
   917 => x"57848080",
   918 => x"81842d76",
   919 => x"80ffffff",
   920 => x"f8065473",
   921 => x"80ffffff",
   922 => x"f82e9438",
   923 => x"fe179fe5",
   924 => x"f408299f",
   925 => x"e5fc0805",
   926 => x"55848080",
   927 => x"9ac50480",
   928 => x"54739fe0",
   929 => x"800c02b4",
   930 => x"050d0402",
   931 => x"e4050d78",
   932 => x"7a71549f",
   933 => x"e5c85355",
   934 => x"55848080",
   935 => x"9a8f2d9f",
   936 => x"e0800881",
   937 => x"ff065372",
   938 => x"802e80fe",
   939 => x"38848080",
   940 => x"a3b45184",
   941 => x"808085ab",
   942 => x"2d9fe5cc",
   943 => x"0883ff05",
   944 => x"892a5780",
   945 => x"70565675",
   946 => x"772580fd",
   947 => x"389fe5d0",
   948 => x"08fe059f",
   949 => x"e5f40829",
   950 => x"9fe5fc08",
   951 => x"11769fe5",
   952 => x"e8080605",
   953 => x"75545253",
   954 => x"8480808e",
   955 => x"a52d9fe0",
   956 => x"8008802e",
   957 => x"80c83881",
   958 => x"15709fe5",
   959 => x"e8080654",
   960 => x"55729438",
   961 => x"9fe5d008",
   962 => x"51848080",
   963 => x"98f92d9f",
   964 => x"e080089f",
   965 => x"e5d00c84",
   966 => x"80148117",
   967 => x"57547676",
   968 => x"24ffaa38",
   969 => x"8480809e",
   970 => x"c9047452",
   971 => x"848080a3",
   972 => x"d0518480",
   973 => x"8081842d",
   974 => x"8480809e",
   975 => x"cb049fe0",
   976 => x"80085384",
   977 => x"80809ecb",
   978 => x"04815372",
   979 => x"9fe0800c",
   980 => x"029c050d",
   981 => x"049fe08c",
   982 => x"08029fe0",
   983 => x"8c0cff3d",
   984 => x"0d800b9f",
   985 => x"e08c08fc",
   986 => x"050c9fe0",
   987 => x"8c088805",
   988 => x"088106ff",
   989 => x"11700970",
   990 => x"9fe08c08",
   991 => x"8c050806",
   992 => x"9fe08c08",
   993 => x"fc050811",
   994 => x"9fe08c08",
   995 => x"fc050c9f",
   996 => x"e08c0888",
   997 => x"0508812a",
   998 => x"9fe08c08",
   999 => x"88050c9f",
  1000 => x"e08c088c",
  1001 => x"0508109f",
  1002 => x"e08c088c",
  1003 => x"050c5151",
  1004 => x"51519fe0",
  1005 => x"8c088805",
  1006 => x"08802e84",
  1007 => x"38ffab39",
  1008 => x"9fe08c08",
  1009 => x"fc050870",
  1010 => x"9fe0800c",
  1011 => x"51833d0d",
  1012 => x"9fe08c0c",
  1013 => x"04000000",
  1014 => x"00ffffff",
  1015 => x"ff00ffff",
  1016 => x"ffff00ff",
  1017 => x"ffffff00",
  1018 => x"436d645f",
  1019 => x"696e6974",
  1020 => x"0a000000",
  1021 => x"496e6974",
  1022 => x"69616c69",
  1023 => x"7a696e67",
  1024 => x"20534420",
  1025 => x"63617264",
  1026 => x"0a000000",
  1027 => x"48756e74",
  1028 => x"696e6720",
  1029 => x"666f7220",
  1030 => x"70617274",
  1031 => x"6974696f",
  1032 => x"6e0a0000",
  1033 => x"4f53445a",
  1034 => x"50553031",
  1035 => x"53595300",
  1036 => x"43616e27",
  1037 => x"74206c6f",
  1038 => x"61642066",
  1039 => x"69726d77",
  1040 => x"6172650a",
  1041 => x"00000000",
  1042 => x"4661696c",
  1043 => x"65642074",
  1044 => x"6f20696e",
  1045 => x"69746961",
  1046 => x"6c697a65",
  1047 => x"20534420",
  1048 => x"63617264",
  1049 => x"0a000000",
  1050 => x"52656164",
  1051 => x"696e6720",
  1052 => x"4d42520a",
  1053 => x"00000000",
  1054 => x"52656164",
  1055 => x"206f6620",
  1056 => x"4d425220",
  1057 => x"6661696c",
  1058 => x"65640a00",
  1059 => x"4d425220",
  1060 => x"73756363",
  1061 => x"65737366",
  1062 => x"756c6c79",
  1063 => x"20726561",
  1064 => x"640a0000",
  1065 => x"46415431",
  1066 => x"36202020",
  1067 => x"00000000",
  1068 => x"46415433",
  1069 => x"32202020",
  1070 => x"00000000",
  1071 => x"50617274",
  1072 => x"6974696f",
  1073 => x"6e636f75",
  1074 => x"6e742025",
  1075 => x"640a0000",
  1076 => x"4e6f2070",
  1077 => x"61727469",
  1078 => x"74696f6e",
  1079 => x"20736967",
  1080 => x"6e617475",
  1081 => x"72652066",
  1082 => x"6f756e64",
  1083 => x"0a000000",
  1084 => x"52656164",
  1085 => x"696e6720",
  1086 => x"626f6f74",
  1087 => x"20736563",
  1088 => x"746f7220",
  1089 => x"25640a00",
  1090 => x"52656164",
  1091 => x"20626f6f",
  1092 => x"74207365",
  1093 => x"63746f72",
  1094 => x"2066726f",
  1095 => x"6d206669",
  1096 => x"72737420",
  1097 => x"70617274",
  1098 => x"6974696f",
  1099 => x"6e0a0000",
  1100 => x"48756e74",
  1101 => x"696e6720",
  1102 => x"666f7220",
  1103 => x"66696c65",
  1104 => x"73797374",
  1105 => x"656d0a00",
  1106 => x"556e7375",
  1107 => x"70706f72",
  1108 => x"74656420",
  1109 => x"70617274",
  1110 => x"6974696f",
  1111 => x"6e207479",
  1112 => x"7065210d",
  1113 => x"00000000",
  1114 => x"52656164",
  1115 => x"696e6720",
  1116 => x"64697265",
  1117 => x"63746f72",
  1118 => x"79207365",
  1119 => x"63746f72",
  1120 => x"2025640a",
  1121 => x"00000000",
  1122 => x"66696c65",
  1123 => x"20222573",
  1124 => x"2220666f",
  1125 => x"756e640d",
  1126 => x"00000000",
  1127 => x"47657446",
  1128 => x"41544c69",
  1129 => x"6e6b2072",
  1130 => x"65747572",
  1131 => x"6e656420",
  1132 => x"25640a00",
  1133 => x"4f70656e",
  1134 => x"65642066",
  1135 => x"696c652c",
  1136 => x"206c6f61",
  1137 => x"64696e67",
  1138 => x"2e2e2e0a",
  1139 => x"00000000",
  1140 => x"43616e27",
  1141 => x"74206f70",
  1142 => x"656e2025",
  1143 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

