-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity DiagROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end DiagROM_ROM;

architecture arch of DiagROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808088",
     1 => x"e8040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90088480",
    10 => x"8088e408",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b848080",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"84808088",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"09810584",
    90 => x"8080889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"84808095",
   162 => x"d0738306",
   163 => x"10100508",
   164 => x"06848080",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"8480808f",
   171 => x"872d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"84808091",
   179 => x"af2d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"80048480",
   279 => x"8088da04",
   280 => x"04000000",
   281 => x"40000460",
   282 => x"84808088",
   283 => x"da0b8480",
   284 => x"8088f404",
   285 => x"02fc050d",
   286 => x"84808095",
   287 => x"e0518480",
   288 => x"80898a2d",
   289 => x"84808089",
   290 => x"840402e0",
   291 => x"050d7958",
   292 => x"77802e90",
   293 => x"38778480",
   294 => x"8095f00c",
   295 => x"800b8480",
   296 => x"8095f80c",
   297 => x"84808095",
   298 => x"f8085271",
   299 => x"82c83884",
   300 => x"808095f0",
   301 => x"08841184",
   302 => x"808095f0",
   303 => x"0c700884",
   304 => x"808095f4",
   305 => x"0c518112",
   306 => x"83068480",
   307 => x"8095f408",
   308 => x"70982c53",
   309 => x"5754800b",
   310 => x"84808095",
   311 => x"f0085355",
   312 => x"70802eaf",
   313 => x"38738480",
   314 => x"8095f80c",
   315 => x"81155573",
   316 => x"81e53871",
   317 => x"84137108",
   318 => x"84808095",
   319 => x"f40c8116",
   320 => x"83068480",
   321 => x"8095f408",
   322 => x"70982c55",
   323 => x"59565353",
   324 => x"70d33871",
   325 => x"84808095",
   326 => x"f00c810b",
   327 => x"82167072",
   328 => x"2a828080",
   329 => x"07595653",
   330 => x"900b86e9",
   331 => x"808423a0",
   332 => x"810b86e9",
   333 => x"80802386",
   334 => x"e9808022",
   335 => x"51800b86",
   336 => x"e9808023",
   337 => x"86e98080",
   338 => x"2252800b",
   339 => x"86e98080",
   340 => x"2386e980",
   341 => x"80227083",
   342 => x"ffff0672",
   343 => x"882a7081",
   344 => x"06515351",
   345 => x"5270802e",
   346 => x"80e03872",
   347 => x"802e81cf",
   348 => x"38718280",
   349 => x"862e0981",
   350 => x"0681a938",
   351 => x"8053fed5",
   352 => x"ca0b86e9",
   353 => x"80802386",
   354 => x"e9808022",
   355 => x"51810b86",
   356 => x"e9808023",
   357 => x"86e98080",
   358 => x"22517286",
   359 => x"e9808023",
   360 => x"86e98080",
   361 => x"22517486",
   362 => x"e9808023",
   363 => x"86e98080",
   364 => x"22517286",
   365 => x"e9808023",
   366 => x"86e98080",
   367 => x"22517286",
   368 => x"e9808023",
   369 => x"86e98080",
   370 => x"2251910b",
   371 => x"86e98084",
   372 => x"23848080",
   373 => x"8aa80475",
   374 => x"882b8480",
   375 => x"8095f40c",
   376 => x"81148306",
   377 => x"84808095",
   378 => x"f4087098",
   379 => x"2c535754",
   380 => x"8480808a",
   381 => x"90048480",
   382 => x"8095f408",
   383 => x"882b8480",
   384 => x"8095f40c",
   385 => x"81128306",
   386 => x"84808095",
   387 => x"f4087098",
   388 => x"2c535754",
   389 => x"800b8480",
   390 => x"8095f008",
   391 => x"53558480",
   392 => x"8089e004",
   393 => x"73848080",
   394 => x"95f80c91",
   395 => x"0b86e980",
   396 => x"8423800b",
   397 => x"84808080",
   398 => x"880c02a0",
   399 => x"050d0476",
   400 => x"722e0981",
   401 => x"06de3871",
   402 => x"1083fe06",
   403 => x"5277802e",
   404 => x"81ee3877",
   405 => x"84808095",
   406 => x"f00c7284",
   407 => x"808095f8",
   408 => x"0c848080",
   409 => x"95f80853",
   410 => x"7281c638",
   411 => x"84808095",
   412 => x"f0088411",
   413 => x"84808095",
   414 => x"f00c7008",
   415 => x"84808095",
   416 => x"f40c5481",
   417 => x"13830684",
   418 => x"808095f8",
   419 => x"0c848080",
   420 => x"95f40870",
   421 => x"982cff14",
   422 => x"54545471",
   423 => x"ff2e80d9",
   424 => x"38848080",
   425 => x"95f00855",
   426 => x"7286e980",
   427 => x"803486e9",
   428 => x"80803351",
   429 => x"72802eae",
   430 => x"38848080",
   431 => x"95f80853",
   432 => x"7280ca38",
   433 => x"74841671",
   434 => x"08848080",
   435 => x"95f40c81",
   436 => x"15830684",
   437 => x"808095f8",
   438 => x"0c848080",
   439 => x"95f40870",
   440 => x"982c5656",
   441 => x"5656ff12",
   442 => x"5271ff2e",
   443 => x"098106ff",
   444 => x"b7387484",
   445 => x"808095f0",
   446 => x"0c910b86",
   447 => x"e9808423",
   448 => x"810b8480",
   449 => x"8080880c",
   450 => x"02a0050d",
   451 => x"0473882b",
   452 => x"84808095",
   453 => x"f40c8113",
   454 => x"83068480",
   455 => x"8095f80c",
   456 => x"84808095",
   457 => x"f4087098",
   458 => x"2c545484",
   459 => x"80808de6",
   460 => x"0475882b",
   461 => x"84808095",
   462 => x"f40c8480",
   463 => x"808d8304",
   464 => x"73848080",
   465 => x"95f80c84",
   466 => x"80808ce1",
   467 => x"0402f005",
   468 => x"0d86e980",
   469 => x"84539073",
   470 => x"2386e980",
   471 => x"80518071",
   472 => x"23702270",
   473 => x"83ffff06",
   474 => x"53548071",
   475 => x"23702254",
   476 => x"80712370",
   477 => x"22519173",
   478 => x"2371882a",
   479 => x"84808080",
   480 => x"880c0290",
   481 => x"050d0484",
   482 => x"80808094",
   483 => x"08028480",
   484 => x"8080940c",
   485 => x"f93d0d80",
   486 => x"0b848080",
   487 => x"809408fc",
   488 => x"050c8480",
   489 => x"80809408",
   490 => x"88050880",
   491 => x"2580c738",
   492 => x"84808080",
   493 => x"94088805",
   494 => x"08308480",
   495 => x"80809408",
   496 => x"88050c80",
   497 => x"0b848080",
   498 => x"809408f4",
   499 => x"050c8480",
   500 => x"80809408",
   501 => x"fc05088c",
   502 => x"38810b84",
   503 => x"80808094",
   504 => x"08f4050c",
   505 => x"84808080",
   506 => x"9408f405",
   507 => x"08848080",
   508 => x"809408fc",
   509 => x"050c8480",
   510 => x"80809408",
   511 => x"8c050880",
   512 => x"2580c738",
   513 => x"84808080",
   514 => x"94088c05",
   515 => x"08308480",
   516 => x"80809408",
   517 => x"8c050c80",
   518 => x"0b848080",
   519 => x"809408f0",
   520 => x"050c8480",
   521 => x"80809408",
   522 => x"fc05088c",
   523 => x"38810b84",
   524 => x"80808094",
   525 => x"08f0050c",
   526 => x"84808080",
   527 => x"9408f005",
   528 => x"08848080",
   529 => x"809408fc",
   530 => x"050c8053",
   531 => x"84808080",
   532 => x"94088c05",
   533 => x"08528480",
   534 => x"80809408",
   535 => x"88050851",
   536 => x"82983f84",
   537 => x"80808088",
   538 => x"08708480",
   539 => x"80809408",
   540 => x"f8050c54",
   541 => x"84808080",
   542 => x"9408fc05",
   543 => x"08802e94",
   544 => x"38848080",
   545 => x"809408f8",
   546 => x"05083084",
   547 => x"80808094",
   548 => x"08f8050c",
   549 => x"84808080",
   550 => x"9408f805",
   551 => x"08708480",
   552 => x"8080880c",
   553 => x"54893d0d",
   554 => x"84808080",
   555 => x"940c0484",
   556 => x"80808094",
   557 => x"08028480",
   558 => x"8080940c",
   559 => x"fb3d0d80",
   560 => x"0b848080",
   561 => x"809408fc",
   562 => x"050c8480",
   563 => x"80809408",
   564 => x"88050880",
   565 => x"259f3884",
   566 => x"80808094",
   567 => x"08880508",
   568 => x"30848080",
   569 => x"80940888",
   570 => x"050c810b",
   571 => x"84808080",
   572 => x"9408fc05",
   573 => x"0c848080",
   574 => x"8094088c",
   575 => x"05088025",
   576 => x"94388480",
   577 => x"80809408",
   578 => x"8c050830",
   579 => x"84808080",
   580 => x"94088c05",
   581 => x"0c815384",
   582 => x"80808094",
   583 => x"088c0508",
   584 => x"52848080",
   585 => x"80940888",
   586 => x"05085180",
   587 => x"cd3f8480",
   588 => x"80808808",
   589 => x"70848080",
   590 => x"809408f8",
   591 => x"050c5484",
   592 => x"80808094",
   593 => x"08fc0508",
   594 => x"802e9438",
   595 => x"84808080",
   596 => x"9408f805",
   597 => x"08308480",
   598 => x"80809408",
   599 => x"f8050c84",
   600 => x"80808094",
   601 => x"08f80508",
   602 => x"70848080",
   603 => x"80880c54",
   604 => x"873d0d84",
   605 => x"80808094",
   606 => x"0c048480",
   607 => x"80809408",
   608 => x"02848080",
   609 => x"80940cfd",
   610 => x"3d0d810b",
   611 => x"84808080",
   612 => x"9408fc05",
   613 => x"0c800b84",
   614 => x"80808094",
   615 => x"08f8050c",
   616 => x"84808080",
   617 => x"94088c05",
   618 => x"08848080",
   619 => x"80940888",
   620 => x"05082780",
   621 => x"c5388480",
   622 => x"80809408",
   623 => x"fc050880",
   624 => x"2eb83880",
   625 => x"0b848080",
   626 => x"8094088c",
   627 => x"050824aa",
   628 => x"38848080",
   629 => x"8094088c",
   630 => x"05081084",
   631 => x"80808094",
   632 => x"088c050c",
   633 => x"84808080",
   634 => x"9408fc05",
   635 => x"08108480",
   636 => x"80809408",
   637 => x"fc050cff",
   638 => x"a7398480",
   639 => x"80809408",
   640 => x"fc050880",
   641 => x"2e80f938",
   642 => x"84808080",
   643 => x"94088c05",
   644 => x"08848080",
   645 => x"80940888",
   646 => x"050826b9",
   647 => x"38848080",
   648 => x"80940888",
   649 => x"05088480",
   650 => x"80809408",
   651 => x"8c050831",
   652 => x"84808080",
   653 => x"94088805",
   654 => x"0c848080",
   655 => x"809408f8",
   656 => x"05088480",
   657 => x"80809408",
   658 => x"fc050807",
   659 => x"84808080",
   660 => x"9408f805",
   661 => x"0c848080",
   662 => x"809408fc",
   663 => x"0508812a",
   664 => x"84808080",
   665 => x"9408fc05",
   666 => x"0c848080",
   667 => x"8094088c",
   668 => x"0508812a",
   669 => x"84808080",
   670 => x"94088c05",
   671 => x"0cfefb39",
   672 => x"84808080",
   673 => x"94089005",
   674 => x"08802e97",
   675 => x"38848080",
   676 => x"80940888",
   677 => x"05087084",
   678 => x"80808094",
   679 => x"08f4050c",
   680 => x"51953984",
   681 => x"80808094",
   682 => x"08f80508",
   683 => x"70848080",
   684 => x"809408f4",
   685 => x"050c5184",
   686 => x"80808094",
   687 => x"08f40508",
   688 => x"84808080",
   689 => x"880c853d",
   690 => x"0d848080",
   691 => x"80940c04",
   692 => x"00ffffff",
   693 => x"ff00ffff",
   694 => x"ffff00ff",
   695 => x"ffffff00",
   696 => x"48656c6c",
   697 => x"6f2c2077",
   698 => x"6f726c64",
   699 => x"210a0064",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

