-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity DiagROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end DiagROM_ROM;

architecture arch of DiagROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"888080ed",
     1 => x"04000000",
     2 => x"00000000",
     3 => x"0b888080",
     4 => x"88080d80",
     5 => x"04888080",
     6 => x"950471fd",
     7 => x"06087283",
     8 => x"06098105",
     9 => x"8205832b",
    10 => x"2a83ffff",
    11 => x"06520471",
    12 => x"fc060872",
    13 => x"83060981",
    14 => x"05830510",
    15 => x"10102a81",
    16 => x"ff065204",
    17 => x"71fc0608",
    18 => x"0b8880a0",
    19 => x"9c738306",
    20 => x"10100508",
    21 => x"067381ff",
    22 => x"06738306",
    23 => x"09810583",
    24 => x"05101010",
    25 => x"2b0772fc",
    26 => x"060c5151",
    27 => x"04028405",
    28 => x"0b888080",
    29 => x"880c8880",
    30 => x"80950b88",
    31 => x"80919404",
    32 => x"0002c405",
    33 => x"0d0280c0",
    34 => x"059fe0e0",
    35 => x"5b568076",
    36 => x"70840558",
    37 => x"08715e5e",
    38 => x"577c7084",
    39 => x"055e0858",
    40 => x"805b7798",
    41 => x"2a78882b",
    42 => x"59547388",
    43 => x"38765e88",
    44 => x"8083cb04",
    45 => x"7b802e81",
    46 => x"ec38805c",
    47 => x"7380e42e",
    48 => x"9f387380",
    49 => x"e4268d38",
    50 => x"7380e32e",
    51 => x"81903888",
    52 => x"8082eb04",
    53 => x"7380f32e",
    54 => x"80ee3888",
    55 => x"8082eb04",
    56 => x"75841771",
    57 => x"087e5c55",
    58 => x"57527280",
    59 => x"258d38ad",
    60 => x"51888090",
    61 => x"c22d7209",
    62 => x"81055372",
    63 => x"802ebb38",
    64 => x"8755729c",
    65 => x"2a73842b",
    66 => x"54527180",
    67 => x"2e833881",
    68 => x"59897225",
    69 => x"8938b712",
    70 => x"52888082",
    71 => x"a104b012",
    72 => x"5278802e",
    73 => x"88387151",
    74 => x"888090c2",
    75 => x"2dff1555",
    76 => x"748025ce",
    77 => x"38888082",
    78 => x"c104b051",
    79 => x"888090c2",
    80 => x"2d805388",
    81 => x"80838104",
    82 => x"75841771",
    83 => x"0870545c",
    84 => x"57528880",
    85 => x"90d62d7b",
    86 => x"53888083",
    87 => x"81047584",
    88 => x"17710856",
    89 => x"57528880",
    90 => x"83b404a5",
    91 => x"51888090",
    92 => x"c22d7351",
    93 => x"888090c2",
    94 => x"2d821757",
    95 => x"888083be",
    96 => x"0472ff14",
    97 => x"54528072",
    98 => x"25b43879",
    99 => x"7081055b",
   100 => x"888080af",
   101 => x"2d705254",
   102 => x"888090c2",
   103 => x"2d811757",
   104 => x"88808381",
   105 => x"0473a52e",
   106 => x"09810688",
   107 => x"38815c88",
   108 => x"8083be04",
   109 => x"73518880",
   110 => x"90c22d81",
   111 => x"1757811b",
   112 => x"5b837b25",
   113 => x"fddc3873",
   114 => x"fdcf387d",
   115 => x"9fe0800c",
   116 => x"02bc050d",
   117 => x"0402f405",
   118 => x"0d747088",
   119 => x"2a83fe80",
   120 => x"06707298",
   121 => x"2a077288",
   122 => x"2b87fc80",
   123 => x"80067398",
   124 => x"2b81f00a",
   125 => x"06717307",
   126 => x"079fe080",
   127 => x"0c565153",
   128 => x"51028c05",
   129 => x"0d0402f8",
   130 => x"050d7388",
   131 => x"2b83fe80",
   132 => x"06028405",
   133 => x"8e058880",
   134 => x"80af2d71",
   135 => x"079fe080",
   136 => x"0c510288",
   137 => x"050d0402",
   138 => x"f8050d73",
   139 => x"70902b71",
   140 => x"902a079f",
   141 => x"e0800c52",
   142 => x"0288050d",
   143 => x"0402f805",
   144 => x"0d735170",
   145 => x"802e8c38",
   146 => x"709fe1a0",
   147 => x"0c800b9f",
   148 => x"e1a80c9f",
   149 => x"e1a80852",
   150 => x"7197389f",
   151 => x"e1a00884",
   152 => x"119fe1a0",
   153 => x"0c70089f",
   154 => x"e1a40c51",
   155 => x"888084fb",
   156 => x"049fe1a4",
   157 => x"08882b9f",
   158 => x"e1a40c81",
   159 => x"1283069f",
   160 => x"e1a80c9f",
   161 => x"e1a40898",
   162 => x"2c9fe080",
   163 => x"0c028805",
   164 => x"0d0402e8",
   165 => x"050d7770",
   166 => x"52568880",
   167 => x"84bd2d9f",
   168 => x"e0800852",
   169 => x"80537180",
   170 => x"2e953881",
   171 => x"13538051",
   172 => x"888084bd",
   173 => x"2d9fe080",
   174 => x"08528880",
   175 => x"85a60482",
   176 => x"13548155",
   177 => x"900b86e9",
   178 => x"808423a0",
   179 => x"810b86e9",
   180 => x"80802386",
   181 => x"e9808022",
   182 => x"52800b86",
   183 => x"e9808023",
   184 => x"86e98080",
   185 => x"2253800b",
   186 => x"86e98080",
   187 => x"2386e980",
   188 => x"80227083",
   189 => x"ffff0673",
   190 => x"882a7081",
   191 => x"06515451",
   192 => x"5371802e",
   193 => x"81a13874",
   194 => x"802e80df",
   195 => x"38728280",
   196 => x"862e0981",
   197 => x"06819038",
   198 => x"8055fed5",
   199 => x"ca0b86e9",
   200 => x"80802386",
   201 => x"e9808022",
   202 => x"52810b86",
   203 => x"e9808023",
   204 => x"86e98080",
   205 => x"22527486",
   206 => x"e9808023",
   207 => x"86e98080",
   208 => x"22527386",
   209 => x"e9808023",
   210 => x"86e98080",
   211 => x"22527486",
   212 => x"e9808023",
   213 => x"86e98080",
   214 => x"22527486",
   215 => x"e9808023",
   216 => x"86e98080",
   217 => x"22528880",
   218 => x"87a70473",
   219 => x"812a8280",
   220 => x"80075272",
   221 => x"722e0981",
   222 => x"06ad3875",
   223 => x"51888084",
   224 => x"bd2d9fe0",
   225 => x"800853ff",
   226 => x"145473ff",
   227 => x"2ea53872",
   228 => x"86e98080",
   229 => x"3486e980",
   230 => x"80335272",
   231 => x"802ee838",
   232 => x"80518880",
   233 => x"86fd0491",
   234 => x"0b86e980",
   235 => x"84238880",
   236 => x"85c40491",
   237 => x"0b86e980",
   238 => x"8423810b",
   239 => x"9fe0800c",
   240 => x"0298050d",
   241 => x"0402f405",
   242 => x"0d86e980",
   243 => x"8052ff72",
   244 => x"34713353",
   245 => x"ff723472",
   246 => x"882b83fe",
   247 => x"80067233",
   248 => x"7081ff06",
   249 => x"515253ff",
   250 => x"72347271",
   251 => x"07882b72",
   252 => x"337081ff",
   253 => x"06515253",
   254 => x"ff723472",
   255 => x"7107882b",
   256 => x"72337081",
   257 => x"ff067207",
   258 => x"9fe0800c",
   259 => x"5253028c",
   260 => x"050d0402",
   261 => x"ec050d76",
   262 => x"78555574",
   263 => x"86e98080",
   264 => x"349fe1ac",
   265 => x"08853873",
   266 => x"892b5473",
   267 => x"982a5372",
   268 => x"86e98080",
   269 => x"3473902a",
   270 => x"537286e9",
   271 => x"80803473",
   272 => x"882a5372",
   273 => x"86e98080",
   274 => x"347386e9",
   275 => x"80803474",
   276 => x"902a5372",
   277 => x"86e98080",
   278 => x"3486e980",
   279 => x"80337081",
   280 => x"ff065153",
   281 => x"82b8bf54",
   282 => x"7281ff2e",
   283 => x"09810699",
   284 => x"38ff0b86",
   285 => x"e9808034",
   286 => x"86e98080",
   287 => x"337081ff",
   288 => x"06ff1656",
   289 => x"515373e0",
   290 => x"38725288",
   291 => x"80a0ac51",
   292 => x"88808181",
   293 => x"2d729fe0",
   294 => x"800c0294",
   295 => x"050d0402",
   296 => x"fc050d81",
   297 => x"c751ff0b",
   298 => x"86e98080",
   299 => x"34ff1151",
   300 => x"708025f2",
   301 => x"38028405",
   302 => x"0d0402f0",
   303 => x"050d8880",
   304 => x"899f2d81",
   305 => x"9c9f5380",
   306 => x"5287fc80",
   307 => x"f7518880",
   308 => x"88932d9f",
   309 => x"e0800854",
   310 => x"9fe08008",
   311 => x"812e0981",
   312 => x"0680e038",
   313 => x"9fe08008",
   314 => x"528880a0",
   315 => x"bc518880",
   316 => x"81812dff",
   317 => x"0b86e980",
   318 => x"8034820a",
   319 => x"52849c80",
   320 => x"e9518880",
   321 => x"88932d9f",
   322 => x"e080089e",
   323 => x"389fe080",
   324 => x"08528880",
   325 => x"a0c85188",
   326 => x"8081812d",
   327 => x"ff0b86e9",
   328 => x"80803473",
   329 => x"5388808a",
   330 => x"d9049fe0",
   331 => x"80085288",
   332 => x"80a0c851",
   333 => x"88808181",
   334 => x"2d888089",
   335 => x"9f2d8880",
   336 => x"8ad2049f",
   337 => x"e0800852",
   338 => x"8880a0bc",
   339 => x"51888081",
   340 => x"812dff13",
   341 => x"5372feef",
   342 => x"38729fe0",
   343 => x"800c0290",
   344 => x"050d0402",
   345 => x"f4050dff",
   346 => x"0b86e980",
   347 => x"80348880",
   348 => x"a0d45188",
   349 => x"8090d62d",
   350 => x"93538052",
   351 => x"87fc80c1",
   352 => x"51888088",
   353 => x"932d9fe0",
   354 => x"80089e38",
   355 => x"9fe08008",
   356 => x"528880a0",
   357 => x"e0518880",
   358 => x"81812dff",
   359 => x"0b86e980",
   360 => x"80348153",
   361 => x"88808bc4",
   362 => x"049fe080",
   363 => x"08528880",
   364 => x"a0e05188",
   365 => x"8081812d",
   366 => x"8880899f",
   367 => x"2dff1353",
   368 => x"72ffb738",
   369 => x"729fe080",
   370 => x"0c028c05",
   371 => x"0d0402f0",
   372 => x"050d8880",
   373 => x"899f2d83",
   374 => x"aa52849c",
   375 => x"80c85188",
   376 => x"8088932d",
   377 => x"9fe08008",
   378 => x"9fe08008",
   379 => x"538880a0",
   380 => x"ec525388",
   381 => x"8081812d",
   382 => x"72812e09",
   383 => x"8106a438",
   384 => x"888087c5",
   385 => x"2d9fe080",
   386 => x"0883ffff",
   387 => x"06537283",
   388 => x"aa2eb238",
   389 => x"9fe08008",
   390 => x"528880a1",
   391 => x"84518880",
   392 => x"81812d88",
   393 => x"808ae32d",
   394 => x"88808cbe",
   395 => x"04815488",
   396 => x"808dea04",
   397 => x"8880a19c",
   398 => x"51888081",
   399 => x"812d8054",
   400 => x"88808dea",
   401 => x"04ff0b86",
   402 => x"e9808034",
   403 => x"b1538880",
   404 => x"89ba2d9f",
   405 => x"e0800880",
   406 => x"2e818038",
   407 => x"805287fc",
   408 => x"80fa5188",
   409 => x"8088932d",
   410 => x"9fe08008",
   411 => x"80de389f",
   412 => x"e0800852",
   413 => x"8880a1b8",
   414 => x"51888081",
   415 => x"812dff0b",
   416 => x"86e98080",
   417 => x"3486e980",
   418 => x"80337081",
   419 => x"ff067054",
   420 => x"8880a1c4",
   421 => x"53515388",
   422 => x"8081812d",
   423 => x"ff0b86e9",
   424 => x"808034ff",
   425 => x"0b86e980",
   426 => x"8034ff0b",
   427 => x"86e98080",
   428 => x"34ff0b86",
   429 => x"e9808034",
   430 => x"72862a70",
   431 => x"81067056",
   432 => x"51537280",
   433 => x"2ea43888",
   434 => x"808cad04",
   435 => x"9fe08008",
   436 => x"528880a1",
   437 => x"b8518880",
   438 => x"81812d72",
   439 => x"822efed4",
   440 => x"38ff1353",
   441 => x"72fee738",
   442 => x"7254739f",
   443 => x"e0800c02",
   444 => x"90050d04",
   445 => x"02f4050d",
   446 => x"810b9fe1",
   447 => x"ac0ca00b",
   448 => x"86e98088",
   449 => x"34830b86",
   450 => x"e9808434",
   451 => x"8880899f",
   452 => x"2d820b86",
   453 => x"e9808434",
   454 => x"87538052",
   455 => x"84d480c0",
   456 => x"51888088",
   457 => x"932d9fe0",
   458 => x"8008812e",
   459 => x"96387282",
   460 => x"2e098106",
   461 => x"88388053",
   462 => x"88808ef3",
   463 => x"04ff1353",
   464 => x"72d83888",
   465 => x"808bce2d",
   466 => x"9fe08008",
   467 => x"9fe1ac0c",
   468 => x"815287fc",
   469 => x"80d05188",
   470 => x"8088932d",
   471 => x"ff0b86e9",
   472 => x"80803483",
   473 => x"0b86e980",
   474 => x"8434ff0b",
   475 => x"86e98080",
   476 => x"34815372",
   477 => x"9fe0800c",
   478 => x"028c050d",
   479 => x"04800b9f",
   480 => x"e0800c04",
   481 => x"02e4050d",
   482 => x"787a5754",
   483 => x"80765474",
   484 => x"538880a1",
   485 => x"d4525788",
   486 => x"8081812d",
   487 => x"ff0b86e9",
   488 => x"80803482",
   489 => x"0b86e980",
   490 => x"8434810b",
   491 => x"86e98088",
   492 => x"34ff0b86",
   493 => x"e9808034",
   494 => x"735287fc",
   495 => x"80d15188",
   496 => x"8088932d",
   497 => x"80dbc6df",
   498 => x"559fe080",
   499 => x"08772e97",
   500 => x"389fe080",
   501 => x"08537352",
   502 => x"8880a1ec",
   503 => x"51888081",
   504 => x"812d8880",
   505 => x"90b804ff",
   506 => x"0b86e980",
   507 => x"803486e9",
   508 => x"80803370",
   509 => x"81ff0651",
   510 => x"547381fe",
   511 => x"2e098106",
   512 => x"a23880ff",
   513 => x"54888087",
   514 => x"c52d9fe0",
   515 => x"80087670",
   516 => x"8405580c",
   517 => x"ff145473",
   518 => x"8025ea38",
   519 => x"81578880",
   520 => x"90aa04ff",
   521 => x"155574ff",
   522 => x"be38ff0b",
   523 => x"86e98080",
   524 => x"34830b86",
   525 => x"e9808434",
   526 => x"769fe080",
   527 => x"0c029c05",
   528 => x"0d0402fc",
   529 => x"050d7270",
   530 => x"86ea8080",
   531 => x"0c9fe080",
   532 => x"0c028405",
   533 => x"0d0402ec",
   534 => x"050d8077",
   535 => x"56547470",
   536 => x"84055608",
   537 => x"51805370",
   538 => x"982a7188",
   539 => x"2b525271",
   540 => x"802e9738",
   541 => x"7186ea80",
   542 => x"800c8114",
   543 => x"81145454",
   544 => x"837325e3",
   545 => x"38888090",
   546 => x"de04739f",
   547 => x"e0800c02",
   548 => x"94050d04",
   549 => x"02f8050d",
   550 => x"8880a28c",
   551 => x"51888090",
   552 => x"d62d8880",
   553 => x"8df42d9f",
   554 => x"e0800880",
   555 => x"2eb33888",
   556 => x"80a2a451",
   557 => x"888090d6",
   558 => x"2d888092",
   559 => x"bd2d8052",
   560 => x"8880a2bc",
   561 => x"5188809d",
   562 => x"d92d9fe0",
   563 => x"8008802e",
   564 => x"86388880",
   565 => x"808c2d88",
   566 => x"80a2c851",
   567 => x"888090d6",
   568 => x"2d8880a2",
   569 => x"e0518880",
   570 => x"90d62d80",
   571 => x"0b9fe080",
   572 => x"0c028805",
   573 => x"0d0402e8",
   574 => x"050d7779",
   575 => x"7b585555",
   576 => x"80537276",
   577 => x"25ab3874",
   578 => x"70810556",
   579 => x"888080af",
   580 => x"2d747081",
   581 => x"05568880",
   582 => x"80af2d52",
   583 => x"5271712e",
   584 => x"88388151",
   585 => x"888092b3",
   586 => x"04811353",
   587 => x"88809282",
   588 => x"04805170",
   589 => x"9fe0800c",
   590 => x"0298050d",
   591 => x"0402d805",
   592 => x"0dff0b9f",
   593 => x"e5d80c80",
   594 => x"0b9fe5ec",
   595 => x"0c8880a3",
   596 => x"80518880",
   597 => x"90d62d9f",
   598 => x"e1c45280",
   599 => x"5188808f",
   600 => x"842d9fe0",
   601 => x"8008549f",
   602 => x"e0800892",
   603 => x"388880a3",
   604 => x"90518880",
   605 => x"90d62d73",
   606 => x"55888099",
   607 => x"d7048880",
   608 => x"a3a45188",
   609 => x"8090d62d",
   610 => x"8056810b",
   611 => x"9fe1b80c",
   612 => x"88538880",
   613 => x"a3bc529f",
   614 => x"e1fa5188",
   615 => x"8091f62d",
   616 => x"9fe08008",
   617 => x"762e0981",
   618 => x"0689389f",
   619 => x"e080089f",
   620 => x"e1b80c88",
   621 => x"538880a3",
   622 => x"c8529fe2",
   623 => x"96518880",
   624 => x"91f62d9f",
   625 => x"e0800889",
   626 => x"389fe080",
   627 => x"089fe1b8",
   628 => x"0c9fe1b8",
   629 => x"08528880",
   630 => x"a3d45188",
   631 => x"8081812d",
   632 => x"9fe1b808",
   633 => x"802e81b1",
   634 => x"389fe58a",
   635 => x"0b888080",
   636 => x"af2d9fe5",
   637 => x"8b0b8880",
   638 => x"80af2d71",
   639 => x"982b7190",
   640 => x"2b079fe5",
   641 => x"8c0b8880",
   642 => x"80af2d70",
   643 => x"882b7207",
   644 => x"9fe58d0b",
   645 => x"888080af",
   646 => x"2d71079f",
   647 => x"e5c20b88",
   648 => x"8080af2d",
   649 => x"9fe5c30b",
   650 => x"888080af",
   651 => x"2d71882b",
   652 => x"07535f54",
   653 => x"525a5657",
   654 => x"557381ab",
   655 => x"aa2e0981",
   656 => x"06923875",
   657 => x"51888083",
   658 => x"d52d9fe0",
   659 => x"80085688",
   660 => x"8094ea04",
   661 => x"7382d4d5",
   662 => x"2e903888",
   663 => x"80a3e851",
   664 => x"888090d6",
   665 => x"2d888096",
   666 => x"d5047552",
   667 => x"8880a488",
   668 => x"51888081",
   669 => x"812d9fe1",
   670 => x"c4527551",
   671 => x"88808f84",
   672 => x"2d9fe080",
   673 => x"08559fe0",
   674 => x"8008802e",
   675 => x"84c93888",
   676 => x"80a4a051",
   677 => x"888090d6",
   678 => x"2d8880a4",
   679 => x"c8518880",
   680 => x"81812d88",
   681 => x"538880a3",
   682 => x"c8529fe2",
   683 => x"96518880",
   684 => x"91f62d9f",
   685 => x"e080088c",
   686 => x"38810b9f",
   687 => x"e5ec0c88",
   688 => x"8095eb04",
   689 => x"88538880",
   690 => x"a3bc529f",
   691 => x"e1fa5188",
   692 => x"8091f62d",
   693 => x"9fe08008",
   694 => x"802e9038",
   695 => x"8880a4e0",
   696 => x"51888081",
   697 => x"812d8880",
   698 => x"96d5049f",
   699 => x"e5c20b88",
   700 => x"8080af2d",
   701 => x"547380d5",
   702 => x"2e098106",
   703 => x"80d7389f",
   704 => x"e5c30b88",
   705 => x"8080af2d",
   706 => x"547381aa",
   707 => x"2e098106",
   708 => x"80c33880",
   709 => x"0b9fe1c4",
   710 => x"0b888080",
   711 => x"af2d5654",
   712 => x"7481e92e",
   713 => x"83388154",
   714 => x"7481eb2e",
   715 => x"8c388055",
   716 => x"73752e09",
   717 => x"8106839f",
   718 => x"389fe1cf",
   719 => x"0b888080",
   720 => x"af2d5574",
   721 => x"90389fe1",
   722 => x"d00b8880",
   723 => x"80af2d54",
   724 => x"73822e88",
   725 => x"38805588",
   726 => x"8099d704",
   727 => x"9fe1d10b",
   728 => x"888080af",
   729 => x"2d709fe5",
   730 => x"f40cff05",
   731 => x"9fe5e80c",
   732 => x"9fe1d20b",
   733 => x"888080af",
   734 => x"2d9fe1d3",
   735 => x"0b888080",
   736 => x"af2d5876",
   737 => x"05778280",
   738 => x"2905709f",
   739 => x"e5dc0c9f",
   740 => x"e1d40b88",
   741 => x"8080af2d",
   742 => x"709fe5d4",
   743 => x"0c9fe5ec",
   744 => x"08595758",
   745 => x"76802e81",
   746 => x"cc388853",
   747 => x"8880a3c8",
   748 => x"529fe296",
   749 => x"51888091",
   750 => x"f62d9fe0",
   751 => x"80088297",
   752 => x"389fe5f4",
   753 => x"0870842b",
   754 => x"9fe5c40c",
   755 => x"709fe5f0",
   756 => x"0c9fe1e9",
   757 => x"0b888080",
   758 => x"af2d9fe1",
   759 => x"e80b8880",
   760 => x"80af2d71",
   761 => x"82802905",
   762 => x"9fe1ea0b",
   763 => x"888080af",
   764 => x"2d708480",
   765 => x"8029129f",
   766 => x"e1eb0b88",
   767 => x"8080af2d",
   768 => x"7081800a",
   769 => x"2912709f",
   770 => x"e1bc0c9f",
   771 => x"e5d40871",
   772 => x"299fe5dc",
   773 => x"0805709f",
   774 => x"e5fc0c9f",
   775 => x"e1f10b88",
   776 => x"8080af2d",
   777 => x"9fe1f00b",
   778 => x"888080af",
   779 => x"2d718280",
   780 => x"29059fe1",
   781 => x"f20b8880",
   782 => x"80af2d70",
   783 => x"84808029",
   784 => x"129fe1f3",
   785 => x"0b888080",
   786 => x"af2d7098",
   787 => x"2b81f00a",
   788 => x"06720570",
   789 => x"9fe1c00c",
   790 => x"fe117e29",
   791 => x"77059fe5",
   792 => x"e40c5259",
   793 => x"5243545e",
   794 => x"51525952",
   795 => x"5d575957",
   796 => x"888099d5",
   797 => x"049fe1d6",
   798 => x"0b888080",
   799 => x"af2d9fe1",
   800 => x"d50b8880",
   801 => x"80af2d71",
   802 => x"82802905",
   803 => x"709fe5c4",
   804 => x"0c70a029",
   805 => x"83ff0570",
   806 => x"892a709f",
   807 => x"e5f00c9f",
   808 => x"e1db0b88",
   809 => x"8080af2d",
   810 => x"9fe1da0b",
   811 => x"888080af",
   812 => x"2d718280",
   813 => x"2905709f",
   814 => x"e1bc0c7b",
   815 => x"71291e70",
   816 => x"9fe5e40c",
   817 => x"7d9fe1c0",
   818 => x"0c73059f",
   819 => x"e5fc0c55",
   820 => x"5e515155",
   821 => x"55815574",
   822 => x"9fe0800c",
   823 => x"02a8050d",
   824 => x"0402ec05",
   825 => x"0d767087",
   826 => x"2c7180ff",
   827 => x"06575553",
   828 => x"9fe5ec08",
   829 => x"8a387288",
   830 => x"2c7381ff",
   831 => x"06565473",
   832 => x"9fe5d808",
   833 => x"2ea3389f",
   834 => x"e1c4529f",
   835 => x"e5dc0814",
   836 => x"5188808f",
   837 => x"842d9fe0",
   838 => x"8008539f",
   839 => x"e0800880",
   840 => x"2e80c538",
   841 => x"739fe5d8",
   842 => x"0c9fe5ec",
   843 => x"08802e9e",
   844 => x"38748429",
   845 => x"9fe1c405",
   846 => x"70085253",
   847 => x"888083d5",
   848 => x"2d9fe080",
   849 => x"08f00a06",
   850 => x"5588809a",
   851 => x"e6047410",
   852 => x"9fe1c405",
   853 => x"70888080",
   854 => x"9a2d5253",
   855 => x"88808486",
   856 => x"2d9fe080",
   857 => x"08557453",
   858 => x"729fe080",
   859 => x"0c029405",
   860 => x"0d0402cc",
   861 => x"050d7e60",
   862 => x"5e5b8056",
   863 => x"ff0b9fe5",
   864 => x"d80c9fe1",
   865 => x"c0089fe5",
   866 => x"e4085657",
   867 => x"9fe5ec08",
   868 => x"762e8d38",
   869 => x"9fe5f408",
   870 => x"842b5988",
   871 => x"809ba704",
   872 => x"9fe5f008",
   873 => x"842b5980",
   874 => x"5a797927",
   875 => x"81d93879",
   876 => x"8f06a017",
   877 => x"5754739f",
   878 => x"38745288",
   879 => x"80a58051",
   880 => x"88808181",
   881 => x"2d9fe1c4",
   882 => x"52745181",
   883 => x"15558880",
   884 => x"8f842d9f",
   885 => x"e1c45680",
   886 => x"76888080",
   887 => x"af2d5558",
   888 => x"73782e83",
   889 => x"38815873",
   890 => x"81e52e81",
   891 => x"92388170",
   892 => x"7906555c",
   893 => x"73802e81",
   894 => x"86388b16",
   895 => x"888080af",
   896 => x"2d980658",
   897 => x"7780f838",
   898 => x"8b537c52",
   899 => x"75518880",
   900 => x"91f62d9f",
   901 => x"e0800880",
   902 => x"e6389c16",
   903 => x"08518880",
   904 => x"83d52d9f",
   905 => x"e0800884",
   906 => x"1c0c9a16",
   907 => x"8880809a",
   908 => x"2d518880",
   909 => x"84862d9f",
   910 => x"e080089f",
   911 => x"e0800855",
   912 => x"559fe5ec",
   913 => x"08802e9d",
   914 => x"38941688",
   915 => x"80809a2d",
   916 => x"51888084",
   917 => x"862d9fe0",
   918 => x"8008902b",
   919 => x"83fff00a",
   920 => x"06701651",
   921 => x"5473881c",
   922 => x"0c777b0c",
   923 => x"7c528880",
   924 => x"a5a05188",
   925 => x"8081812d",
   926 => x"7b548880",
   927 => x"9dcf0481",
   928 => x"1a5a8880",
   929 => x"9ba9049f",
   930 => x"e5ec0880",
   931 => x"2ebf3876",
   932 => x"51888099",
   933 => x"e12d9fe0",
   934 => x"80089fe0",
   935 => x"80085388",
   936 => x"80a5b452",
   937 => x"57888081",
   938 => x"812d7680",
   939 => x"fffffff8",
   940 => x"06547380",
   941 => x"fffffff8",
   942 => x"2e9338fe",
   943 => x"179fe5f4",
   944 => x"08299fe5",
   945 => x"fc080555",
   946 => x"88809ba7",
   947 => x"04805473",
   948 => x"9fe0800c",
   949 => x"02b4050d",
   950 => x"0402e405",
   951 => x"0d787a71",
   952 => x"549fe5c8",
   953 => x"53555588",
   954 => x"809af22d",
   955 => x"9fe08008",
   956 => x"81ff0653",
   957 => x"72802e80",
   958 => x"f9388880",
   959 => x"a5cc5188",
   960 => x"8090d62d",
   961 => x"9fe5cc08",
   962 => x"83ff0589",
   963 => x"2a578070",
   964 => x"56567577",
   965 => x"2580f638",
   966 => x"9fe5d008",
   967 => x"fe059fe5",
   968 => x"f408299f",
   969 => x"e5fc0811",
   970 => x"769fe5e8",
   971 => x"08060575",
   972 => x"54525388",
   973 => x"808f842d",
   974 => x"9fe08008",
   975 => x"802e80c3",
   976 => x"38811570",
   977 => x"9fe5e808",
   978 => x"06545572",
   979 => x"93389fe5",
   980 => x"d0085188",
   981 => x"8099e12d",
   982 => x"9fe08008",
   983 => x"9fe5d00c",
   984 => x"84801481",
   985 => x"17575476",
   986 => x"7624ffac",
   987 => x"3888809f",
   988 => x"8d047452",
   989 => x"8880a5e8",
   990 => x"51888081",
   991 => x"812d8880",
   992 => x"9f8f049f",
   993 => x"e0800853",
   994 => x"88809f8f",
   995 => x"04815372",
   996 => x"9fe0800c",
   997 => x"029c050d",
   998 => x"049fe08c",
   999 => x"08029fe0",
  1000 => x"8c0cff3d",
  1001 => x"0d800b9f",
  1002 => x"e08c08fc",
  1003 => x"050c9fe0",
  1004 => x"8c088805",
  1005 => x"088106ff",
  1006 => x"11700970",
  1007 => x"9fe08c08",
  1008 => x"8c050806",
  1009 => x"9fe08c08",
  1010 => x"fc050811",
  1011 => x"9fe08c08",
  1012 => x"fc050c9f",
  1013 => x"e08c0888",
  1014 => x"0508812a",
  1015 => x"9fe08c08",
  1016 => x"88050c9f",
  1017 => x"e08c088c",
  1018 => x"0508109f",
  1019 => x"e08c088c",
  1020 => x"050c5151",
  1021 => x"51519fe0",
  1022 => x"8c088805",
  1023 => x"08802e84",
  1024 => x"38ffab39",
  1025 => x"9fe08c08",
  1026 => x"fc050870",
  1027 => x"9fe0800c",
  1028 => x"51833d0d",
  1029 => x"9fe08c0c",
  1030 => x"04000000",
  1031 => x"00ffffff",
  1032 => x"ff00ffff",
  1033 => x"ffff00ff",
  1034 => x"ffffff00",
  1035 => x"476f7420",
  1036 => x"72657375",
  1037 => x"6c742025",
  1038 => x"64200a00",
  1039 => x"434d4435",
  1040 => x"35202564",
  1041 => x"0a000000",
  1042 => x"434d4434",
  1043 => x"31202564",
  1044 => x"0a000000",
  1045 => x"436d645f",
  1046 => x"696e6974",
  1047 => x"0a000000",
  1048 => x"696e6974",
  1049 => x"2025640a",
  1050 => x"20200000",
  1051 => x"636d645f",
  1052 => x"434d4438",
  1053 => x"20726573",
  1054 => x"706f6e73",
  1055 => x"653a2025",
  1056 => x"640a0000",
  1057 => x"434d4438",
  1058 => x"5f342072",
  1059 => x"6573706f",
  1060 => x"6e73653a",
  1061 => x"2025640a",
  1062 => x"00000000",
  1063 => x"53444843",
  1064 => x"20496e69",
  1065 => x"7469616c",
  1066 => x"697a6174",
  1067 => x"696f6e20",
  1068 => x"6572726f",
  1069 => x"72210a00",
  1070 => x"434d4435",
  1071 => x"38202564",
  1072 => x"0a202000",
  1073 => x"434d4435",
  1074 => x"385f3220",
  1075 => x"25640a20",
  1076 => x"20000000",
  1077 => x"73645f72",
  1078 => x"6561645f",
  1079 => x"73656374",
  1080 => x"6f722025",
  1081 => x"642c2025",
  1082 => x"640a0000",
  1083 => x"52656164",
  1084 => x"20636f6d",
  1085 => x"6d616e64",
  1086 => x"20666169",
  1087 => x"6c656420",
  1088 => x"61742025",
  1089 => x"64202825",
  1090 => x"64290a00",
  1091 => x"496e6974",
  1092 => x"69616c69",
  1093 => x"7a696e67",
  1094 => x"20534420",
  1095 => x"63617264",
  1096 => x"0a000000",
  1097 => x"48756e74",
  1098 => x"696e6720",
  1099 => x"666f7220",
  1100 => x"70617274",
  1101 => x"6974696f",
  1102 => x"6e0a0000",
  1103 => x"4f53445a",
  1104 => x"50553031",
  1105 => x"53595300",
  1106 => x"43616e27",
  1107 => x"74206c6f",
  1108 => x"61642066",
  1109 => x"69726d77",
  1110 => x"6172650a",
  1111 => x"00000000",
  1112 => x"4661696c",
  1113 => x"65642074",
  1114 => x"6f20696e",
  1115 => x"69746961",
  1116 => x"6c697a65",
  1117 => x"20534420",
  1118 => x"63617264",
  1119 => x"0a000000",
  1120 => x"52656164",
  1121 => x"696e6720",
  1122 => x"4d42520a",
  1123 => x"00000000",
  1124 => x"52656164",
  1125 => x"206f6620",
  1126 => x"4d425220",
  1127 => x"6661696c",
  1128 => x"65640a00",
  1129 => x"4d425220",
  1130 => x"73756363",
  1131 => x"65737366",
  1132 => x"756c6c79",
  1133 => x"20726561",
  1134 => x"640a0000",
  1135 => x"46415431",
  1136 => x"36202020",
  1137 => x"00000000",
  1138 => x"46415433",
  1139 => x"32202020",
  1140 => x"00000000",
  1141 => x"50617274",
  1142 => x"6974696f",
  1143 => x"6e636f75",
  1144 => x"6e742025",
  1145 => x"640a0000",
  1146 => x"4e6f2070",
  1147 => x"61727469",
  1148 => x"74696f6e",
  1149 => x"20736967",
  1150 => x"6e617475",
  1151 => x"72652066",
  1152 => x"6f756e64",
  1153 => x"0a000000",
  1154 => x"52656164",
  1155 => x"696e6720",
  1156 => x"626f6f74",
  1157 => x"20736563",
  1158 => x"746f7220",
  1159 => x"25640a00",
  1160 => x"52656164",
  1161 => x"20626f6f",
  1162 => x"74207365",
  1163 => x"63746f72",
  1164 => x"2066726f",
  1165 => x"6d206669",
  1166 => x"72737420",
  1167 => x"70617274",
  1168 => x"6974696f",
  1169 => x"6e0a0000",
  1170 => x"48756e74",
  1171 => x"696e6720",
  1172 => x"666f7220",
  1173 => x"66696c65",
  1174 => x"73797374",
  1175 => x"656d0a00",
  1176 => x"556e7375",
  1177 => x"70706f72",
  1178 => x"74656420",
  1179 => x"70617274",
  1180 => x"6974696f",
  1181 => x"6e207479",
  1182 => x"7065210d",
  1183 => x"00000000",
  1184 => x"52656164",
  1185 => x"696e6720",
  1186 => x"64697265",
  1187 => x"63746f72",
  1188 => x"79207365",
  1189 => x"63746f72",
  1190 => x"2025640a",
  1191 => x"00000000",
  1192 => x"66696c65",
  1193 => x"20222573",
  1194 => x"2220666f",
  1195 => x"756e640d",
  1196 => x"00000000",
  1197 => x"47657446",
  1198 => x"41544c69",
  1199 => x"6e6b2072",
  1200 => x"65747572",
  1201 => x"6e656420",
  1202 => x"25640a00",
  1203 => x"4f70656e",
  1204 => x"65642066",
  1205 => x"696c652c",
  1206 => x"206c6f61",
  1207 => x"64696e67",
  1208 => x"2e2e2e0a",
  1209 => x"00000000",
  1210 => x"43616e27",
  1211 => x"74206f70",
  1212 => x"656e2025",
  1213 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

