-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity DiagROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end DiagROM_ROM;

architecture arch of DiagROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ed040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"880d8004",
     5 => x"84808080",
     6 => x"940471fd",
     7 => x"06087283",
     8 => x"06098105",
     9 => x"8205832b",
    10 => x"2a83ffff",
    11 => x"06520471",
    12 => x"fc060872",
    13 => x"83060981",
    14 => x"05830510",
    15 => x"10102a81",
    16 => x"ff065204",
    17 => x"71fc0608",
    18 => x"848080ac",
    19 => x"d0738306",
    20 => x"10100508",
    21 => x"067381ff",
    22 => x"06738306",
    23 => x"09810583",
    24 => x"05101010",
    25 => x"2b0772fc",
    26 => x"060c5151",
    27 => x"04028405",
    28 => x"84808080",
    29 => x"880c8480",
    30 => x"8080940b",
    31 => x"8480809b",
    32 => x"c8040000",
    33 => x"02c4050d",
    34 => x"0280c005",
    35 => x"83ffe0e0",
    36 => x"5b568076",
    37 => x"70840558",
    38 => x"08715e5e",
    39 => x"577c7084",
    40 => x"055e0858",
    41 => x"805b7798",
    42 => x"2a78882b",
    43 => x"59547389",
    44 => x"38765e84",
    45 => x"808083e3",
    46 => x"047b802e",
    47 => x"81fd3880",
    48 => x"5c7380e4",
    49 => x"2ea13873",
    50 => x"80e4268e",
    51 => x"387380e3",
    52 => x"2e819a38",
    53 => x"84808082",
    54 => x"fb047380",
    55 => x"f32e80f5",
    56 => x"38848080",
    57 => x"82fb0475",
    58 => x"84177108",
    59 => x"7e5c5557",
    60 => x"52728025",
    61 => x"8e38ad51",
    62 => x"8480809b",
    63 => x"b92d7209",
    64 => x"81055372",
    65 => x"802ebe38",
    66 => x"8755729c",
    67 => x"2a73842b",
    68 => x"54527180",
    69 => x"2e833881",
    70 => x"59897225",
    71 => x"8a38b712",
    72 => x"52848080",
    73 => x"82aa04b0",
    74 => x"12527880",
    75 => x"2e893871",
    76 => x"51848080",
    77 => x"9bb92dff",
    78 => x"15557480",
    79 => x"25cc3884",
    80 => x"808082cd",
    81 => x"04b05184",
    82 => x"80809bb9",
    83 => x"2d805384",
    84 => x"80808394",
    85 => x"04758417",
    86 => x"71087054",
    87 => x"5c575284",
    88 => x"808086dc",
    89 => x"2d7b5384",
    90 => x"80808394",
    91 => x"04758417",
    92 => x"71085657",
    93 => x"52848080",
    94 => x"83cb04a5",
    95 => x"51848080",
    96 => x"9bb92d73",
    97 => x"51848080",
    98 => x"9bb92d82",
    99 => x"17578480",
   100 => x"8083d604",
   101 => x"72ff1454",
   102 => x"52807225",
   103 => x"b9387970",
   104 => x"81055b84",
   105 => x"808080af",
   106 => x"2d705254",
   107 => x"8480809b",
   108 => x"b92d8117",
   109 => x"57848080",
   110 => x"83940473",
   111 => x"a52e0981",
   112 => x"06893881",
   113 => x"5c848080",
   114 => x"83d60473",
   115 => x"51848080",
   116 => x"9bb92d81",
   117 => x"1757811b",
   118 => x"5b837b25",
   119 => x"fdc83873",
   120 => x"fdbb387d",
   121 => x"83ffe080",
   122 => x"0c02bc05",
   123 => x"0d0402f4",
   124 => x"050d7470",
   125 => x"882a83fe",
   126 => x"80067072",
   127 => x"982a0772",
   128 => x"882b87fc",
   129 => x"80800673",
   130 => x"982b81f0",
   131 => x"0a067173",
   132 => x"070783ff",
   133 => x"e0800c56",
   134 => x"51535102",
   135 => x"8c050d04",
   136 => x"02f8050d",
   137 => x"028e0584",
   138 => x"808080af",
   139 => x"2d74982b",
   140 => x"71902b07",
   141 => x"70902c83",
   142 => x"ffe0800c",
   143 => x"52520288",
   144 => x"050d0402",
   145 => x"f8050d73",
   146 => x"70902b71",
   147 => x"902a0783",
   148 => x"ffe0800c",
   149 => x"52028805",
   150 => x"0d0483ff",
   151 => x"e08c0802",
   152 => x"83ffe08c",
   153 => x"0c803d0d",
   154 => x"83ffe08c",
   155 => x"08880508",
   156 => x"802e9538",
   157 => x"83ffe08c",
   158 => x"08880508",
   159 => x"83ffe1a0",
   160 => x"0c800b83",
   161 => x"ffe1a80c",
   162 => x"83ffe1a8",
   163 => x"089c3883",
   164 => x"ffe1a008",
   165 => x"83ffe1a0",
   166 => x"08840583",
   167 => x"ffe1a00c",
   168 => x"700883ff",
   169 => x"e1a40c51",
   170 => x"8d3983ff",
   171 => x"e1a40888",
   172 => x"2b83ffe1",
   173 => x"a40c83ff",
   174 => x"e1a80881",
   175 => x"05708306",
   176 => x"83ffe1a8",
   177 => x"0c83ffe1",
   178 => x"a408982c",
   179 => x"7083ffe0",
   180 => x"800c5151",
   181 => x"823d0d83",
   182 => x"ffe08c0c",
   183 => x"0483ffe0",
   184 => x"8c080283",
   185 => x"ffe08c0c",
   186 => x"fd3d0d83",
   187 => x"ffe08c08",
   188 => x"88050851",
   189 => x"fee43f83",
   190 => x"ffe08008",
   191 => x"7083ffe0",
   192 => x"8c08fc05",
   193 => x"0c52800b",
   194 => x"83ffe08c",
   195 => x"08f8050c",
   196 => x"83ffe08c",
   197 => x"08fc0508",
   198 => x"802ea938",
   199 => x"83ffe08c",
   200 => x"08f80508",
   201 => x"810583ff",
   202 => x"e08c08f8",
   203 => x"050c8051",
   204 => x"fea83f83",
   205 => x"ffe08008",
   206 => x"7083ffe0",
   207 => x"8c08fc05",
   208 => x"0c52cd39",
   209 => x"83ffe08c",
   210 => x"08f80508",
   211 => x"7083ffe0",
   212 => x"800c5285",
   213 => x"3d0d83ff",
   214 => x"e08c0c04",
   215 => x"83ffe08c",
   216 => x"080283ff",
   217 => x"e08c0cf7",
   218 => x"3d0d83ff",
   219 => x"e08c0888",
   220 => x"050883ff",
   221 => x"e08c08e8",
   222 => x"050c83ff",
   223 => x"e08c0888",
   224 => x"050851fe",
   225 => x"d83f83ff",
   226 => x"e0800882",
   227 => x"1183ffe0",
   228 => x"8c08e405",
   229 => x"0c52810b",
   230 => x"83ffe08c",
   231 => x"08ec050c",
   232 => x"900b86e9",
   233 => x"808423a0",
   234 => x"810b86e9",
   235 => x"80802386",
   236 => x"e9808022",
   237 => x"7083ffff",
   238 => x"0683ffe0",
   239 => x"8c08fc05",
   240 => x"0c52800b",
   241 => x"86e98080",
   242 => x"2386e980",
   243 => x"80225280",
   244 => x"0b86e980",
   245 => x"802386e9",
   246 => x"80802270",
   247 => x"83ffff06",
   248 => x"83ffe08c",
   249 => x"08f4050c",
   250 => x"83ffe08c",
   251 => x"08fc0508",
   252 => x"882a7081",
   253 => x"06515152",
   254 => x"71802e82",
   255 => x"b73883ff",
   256 => x"e08c08ec",
   257 => x"0508802e",
   258 => x"80f83883",
   259 => x"ffe08c08",
   260 => x"f4050882",
   261 => x"80862e09",
   262 => x"81068298",
   263 => x"38800b83",
   264 => x"ffe08c08",
   265 => x"ec050cfe",
   266 => x"d5ca0b86",
   267 => x"e9808023",
   268 => x"86e98080",
   269 => x"2252810b",
   270 => x"86e98080",
   271 => x"2386e980",
   272 => x"80225280",
   273 => x"0b86e980",
   274 => x"802386e9",
   275 => x"80802283",
   276 => x"ffe08c08",
   277 => x"e4050851",
   278 => x"527186e9",
   279 => x"80802386",
   280 => x"e9808022",
   281 => x"52800b86",
   282 => x"e9808023",
   283 => x"86e98080",
   284 => x"2252800b",
   285 => x"86e98080",
   286 => x"2386e980",
   287 => x"80225281",
   288 => x"b33983ff",
   289 => x"e08c08e4",
   290 => x"0508812a",
   291 => x"70828080",
   292 => x"07515271",
   293 => x"83ffe08c",
   294 => x"08f40508",
   295 => x"2e098106",
   296 => x"81923883",
   297 => x"ffe08c08",
   298 => x"f0050810",
   299 => x"83ffe08c",
   300 => x"08e4050c",
   301 => x"83ffe08c",
   302 => x"08880508",
   303 => x"51fb9b3f",
   304 => x"83ffe080",
   305 => x"0883ffe0",
   306 => x"8c08f005",
   307 => x"0c83ffe0",
   308 => x"8c08e405",
   309 => x"08ff0583",
   310 => x"ffe08c08",
   311 => x"e4050c83",
   312 => x"ffe08c08",
   313 => x"e40508ff",
   314 => x"2eb73883",
   315 => x"ffe08c08",
   316 => x"f0050852",
   317 => x"7186e980",
   318 => x"803486e9",
   319 => x"80803352",
   320 => x"83ffe08c",
   321 => x"08f00508",
   322 => x"802ec238",
   323 => x"8051faca",
   324 => x"3f83ffe0",
   325 => x"800883ff",
   326 => x"e08c08f0",
   327 => x"050cffad",
   328 => x"39910b86",
   329 => x"e9808423",
   330 => x"810b83ff",
   331 => x"e08c08e0",
   332 => x"050c8b39",
   333 => x"910b86e9",
   334 => x"808423fc",
   335 => x"e33983ff",
   336 => x"e08c08e0",
   337 => x"050883ff",
   338 => x"e0800c8b",
   339 => x"3d0d83ff",
   340 => x"e08c0c04",
   341 => x"83ffe08c",
   342 => x"080283ff",
   343 => x"e08c0cfe",
   344 => x"3d0d800b",
   345 => x"83ffe08c",
   346 => x"08fc050c",
   347 => x"81ff0b86",
   348 => x"e9808023",
   349 => x"86e98080",
   350 => x"227083ff",
   351 => x"ff067081",
   352 => x"ff0683ff",
   353 => x"e08c08fc",
   354 => x"050c5151",
   355 => x"81ff0b86",
   356 => x"e9808023",
   357 => x"83ffe08c",
   358 => x"08fc0508",
   359 => x"882b5286",
   360 => x"e9808022",
   361 => x"7083ffff",
   362 => x"067081ff",
   363 => x"06707507",
   364 => x"83ffe08c",
   365 => x"08fc050c",
   366 => x"51515181",
   367 => x"ff0b86e9",
   368 => x"80802383",
   369 => x"ffe08c08",
   370 => x"fc050888",
   371 => x"2b5286e9",
   372 => x"80802270",
   373 => x"83ffff06",
   374 => x"7081ff06",
   375 => x"70750783",
   376 => x"ffe08c08",
   377 => x"fc050c51",
   378 => x"515181ff",
   379 => x"0b86e980",
   380 => x"802383ff",
   381 => x"e08c08fc",
   382 => x"0508882b",
   383 => x"5286e980",
   384 => x"80227083",
   385 => x"ffff0670",
   386 => x"81ff0670",
   387 => x"750783ff",
   388 => x"e08c08fc",
   389 => x"050c83ff",
   390 => x"e08c08fc",
   391 => x"05087083",
   392 => x"ffe0800c",
   393 => x"51515151",
   394 => x"843d0d83",
   395 => x"ffe08c0c",
   396 => x"0483ffe0",
   397 => x"8c080283",
   398 => x"ffe08c0c",
   399 => x"fe3d0d81",
   400 => x"ff0b83ff",
   401 => x"e08c08f8",
   402 => x"050c83ff",
   403 => x"e08c0888",
   404 => x"05087081",
   405 => x"ff065151",
   406 => x"7086e980",
   407 => x"802383ff",
   408 => x"e1ac0893",
   409 => x"3883ffe0",
   410 => x"8c088c05",
   411 => x"08892b83",
   412 => x"ffe08c08",
   413 => x"8c050c83",
   414 => x"ffe08c08",
   415 => x"8c050898",
   416 => x"2a7081ff",
   417 => x"06515170",
   418 => x"86e98080",
   419 => x"2383ffe0",
   420 => x"8c088c05",
   421 => x"08902a70",
   422 => x"81ff0651",
   423 => x"517086e9",
   424 => x"80802383",
   425 => x"ffe08c08",
   426 => x"8c050888",
   427 => x"2a7081ff",
   428 => x"06515170",
   429 => x"86e98080",
   430 => x"2383ffe0",
   431 => x"8c088c05",
   432 => x"087081ff",
   433 => x"06515170",
   434 => x"86e98080",
   435 => x"2383ffe0",
   436 => x"8c088805",
   437 => x"08902a70",
   438 => x"81ff0651",
   439 => x"517086e9",
   440 => x"80802382",
   441 => x"b8c00b83",
   442 => x"ffe08c08",
   443 => x"fc050c86",
   444 => x"e9808022",
   445 => x"7083ffff",
   446 => x"067081ff",
   447 => x"0683ffe0",
   448 => x"8c08f805",
   449 => x"0c515183",
   450 => x"ffe08c08",
   451 => x"fc0508ff",
   452 => x"0583ffe0",
   453 => x"8c08fc05",
   454 => x"0c83ffe0",
   455 => x"8c08fc05",
   456 => x"08802eb4",
   457 => x"3883ffe0",
   458 => x"8c08f805",
   459 => x"0881ff2e",
   460 => x"098106a4",
   461 => x"3881ff0b",
   462 => x"86e98080",
   463 => x"2386e980",
   464 => x"80227083",
   465 => x"ffff0670",
   466 => x"81ff0683",
   467 => x"ffe08c08",
   468 => x"f8050c51",
   469 => x"51ffb039",
   470 => x"83ffe08c",
   471 => x"08f80508",
   472 => x"7083ffe0",
   473 => x"800c5184",
   474 => x"3d0d83ff",
   475 => x"e08c0c04",
   476 => x"83ffe08c",
   477 => x"080283ff",
   478 => x"e08c0c80",
   479 => x"3d0d800b",
   480 => x"83ffe08c",
   481 => x"08fc050c",
   482 => x"83ffe08c",
   483 => x"08fc0508",
   484 => x"81c7249d",
   485 => x"3881ff0b",
   486 => x"86e98080",
   487 => x"2383ffe0",
   488 => x"8c08fc05",
   489 => x"08810583",
   490 => x"ffe08c08",
   491 => x"fc050cd8",
   492 => x"39823d0d",
   493 => x"83ffe08c",
   494 => x"0c0483ff",
   495 => x"e08c0802",
   496 => x"83ffe08c",
   497 => x"0cfb3d0d",
   498 => x"819ca00b",
   499 => x"83ffe08c",
   500 => x"08fc050c",
   501 => x"ff9a3f83",
   502 => x"ffe08c08",
   503 => x"fc0508ff",
   504 => x"0583ffe0",
   505 => x"8c08fc05",
   506 => x"0c83ffe0",
   507 => x"8c08fc05",
   508 => x"08802e80",
   509 => x"f0388052",
   510 => x"87fc80f7",
   511 => x"51fcb23f",
   512 => x"83ffe080",
   513 => x"087083ff",
   514 => x"e08c08f8",
   515 => x"050c5383",
   516 => x"ffe08c08",
   517 => x"f8050881",
   518 => x"2e098106",
   519 => x"ffb93881",
   520 => x"ff0b86e9",
   521 => x"80802382",
   522 => x"0a52849c",
   523 => x"80e951fc",
   524 => x"803f83ff",
   525 => x"e0800870",
   526 => x"83ffe08c",
   527 => x"08f8050c",
   528 => x"5383ffe0",
   529 => x"8c08f805",
   530 => x"08953881",
   531 => x"ff0b86e9",
   532 => x"80802381",
   533 => x"0b83ffe0",
   534 => x"8c08f405",
   535 => x"0c9139fe",
   536 => x"8f3ffef3",
   537 => x"39800b83",
   538 => x"ffe08c08",
   539 => x"f4050c83",
   540 => x"ffe08c08",
   541 => x"f4050883",
   542 => x"ffe0800c",
   543 => x"873d0d83",
   544 => x"ffe08c0c",
   545 => x"0483ffe0",
   546 => x"8c080283",
   547 => x"ffe08c0c",
   548 => x"fb3d0d94",
   549 => x"0b83ffe0",
   550 => x"8c08fc05",
   551 => x"0c81ff0b",
   552 => x"86e98080",
   553 => x"23848080",
   554 => x"ace051f5",
   555 => x"af3f83ff",
   556 => x"e08c08fc",
   557 => x"0508ff05",
   558 => x"83ffe08c",
   559 => x"08fc050c",
   560 => x"83ffe08c",
   561 => x"08fc0508",
   562 => x"802ebe38",
   563 => x"805287fc",
   564 => x"80c151fa",
   565 => x"dc3f83ff",
   566 => x"e0800870",
   567 => x"83ffe08c",
   568 => x"08f8050c",
   569 => x"5383ffe0",
   570 => x"8c08f805",
   571 => x"08953881",
   572 => x"ff0b86e9",
   573 => x"80802381",
   574 => x"0b83ffe0",
   575 => x"8c08f405",
   576 => x"0c9139fc",
   577 => x"eb3fffa6",
   578 => x"39800b83",
   579 => x"ffe08c08",
   580 => x"f4050c83",
   581 => x"ffe08c08",
   582 => x"f4050883",
   583 => x"ffe0800c",
   584 => x"873d0d83",
   585 => x"ffe08c0c",
   586 => x"0483ffe0",
   587 => x"8c080283",
   588 => x"ffe08c0c",
   589 => x"fb3d0dfc",
   590 => x"b73f83aa",
   591 => x"52849c80",
   592 => x"c851f9ed",
   593 => x"3f83ffe0",
   594 => x"80087083",
   595 => x"ffe08c08",
   596 => x"f8050c83",
   597 => x"ffe08c08",
   598 => x"f8050853",
   599 => x"848080ac",
   600 => x"ec5253ee",
   601 => x"9f3f83ff",
   602 => x"e08c08f8",
   603 => x"0508812e",
   604 => x"9138fe91",
   605 => x"3f800b83",
   606 => x"ffe08c08",
   607 => x"f4050c82",
   608 => x"ff39f7d0",
   609 => x"3f83ffe0",
   610 => x"80087083",
   611 => x"ffe08c08",
   612 => x"f8050c83",
   613 => x"ffe08c08",
   614 => x"f8050883",
   615 => x"ffff0651",
   616 => x"537283aa",
   617 => x"2ea33883",
   618 => x"ffe08c08",
   619 => x"f8050852",
   620 => x"848080ad",
   621 => x"8451edcc",
   622 => x"3ffdca3f",
   623 => x"800b83ff",
   624 => x"e08c08f4",
   625 => x"050c82b8",
   626 => x"3981ff0b",
   627 => x"86e98080",
   628 => x"23b20b83",
   629 => x"ffe08c08",
   630 => x"fc050c83",
   631 => x"ffe08c08",
   632 => x"fc0508ff",
   633 => x"0583ffe0",
   634 => x"8c08fc05",
   635 => x"0c83ffe0",
   636 => x"8c08fc05",
   637 => x"08802e81",
   638 => x"fd38fbbe",
   639 => x"3f83ffe0",
   640 => x"80085372",
   641 => x"802e81c9",
   642 => x"38805287",
   643 => x"fc80fa51",
   644 => x"f89f3f83",
   645 => x"ffe08008",
   646 => x"7083ffe0",
   647 => x"8c08f805",
   648 => x"0c5383ff",
   649 => x"e08c08f8",
   650 => x"05088193",
   651 => x"3883ffe0",
   652 => x"8c08f805",
   653 => x"08528480",
   654 => x"80ad9c51",
   655 => x"ecc63f81",
   656 => x"ff0b86e9",
   657 => x"80802386",
   658 => x"e9808022",
   659 => x"7083ffff",
   660 => x"067081ff",
   661 => x"0683ffe0",
   662 => x"8c08f805",
   663 => x"0c83ffe0",
   664 => x"8c08f805",
   665 => x"08548480",
   666 => x"80ada853",
   667 => x"5153ec94",
   668 => x"3f81ff0b",
   669 => x"86e98080",
   670 => x"2381ff0b",
   671 => x"86e98080",
   672 => x"2381ff0b",
   673 => x"86e98080",
   674 => x"2381ff0b",
   675 => x"86e98080",
   676 => x"2383ffe0",
   677 => x"8c08f805",
   678 => x"08862a70",
   679 => x"81065153",
   680 => x"72802e8e",
   681 => x"38810b83",
   682 => x"ffe08c08",
   683 => x"f4050c80",
   684 => x"cf39800b",
   685 => x"83ffe08c",
   686 => x"08f4050c",
   687 => x"80c23983",
   688 => x"ffe08c08",
   689 => x"f8050852",
   690 => x"848080ad",
   691 => x"9c51ebb4",
   692 => x"3f83ffe0",
   693 => x"8c08fc05",
   694 => x"08822e09",
   695 => x"8106fdfb",
   696 => x"38848080",
   697 => x"adb851eb",
   698 => x"9b3f800b",
   699 => x"83ffe08c",
   700 => x"08f4050c",
   701 => x"8b39800b",
   702 => x"83ffe08c",
   703 => x"08f4050c",
   704 => x"83ffe08c",
   705 => x"08f40508",
   706 => x"83ffe080",
   707 => x"0c873d0d",
   708 => x"83ffe08c",
   709 => x"0c0483ff",
   710 => x"e08c0802",
   711 => x"83ffe08c",
   712 => x"0cfb3d0d",
   713 => x"810b83ff",
   714 => x"e1ac0ca0",
   715 => x"0b86e980",
   716 => x"8823830b",
   717 => x"86e98084",
   718 => x"23f8b53f",
   719 => x"820b86e9",
   720 => x"80842388",
   721 => x"0b83ffe0",
   722 => x"8c08fc05",
   723 => x"0c83ffe0",
   724 => x"8c08fc05",
   725 => x"08ff0583",
   726 => x"ffe08c08",
   727 => x"fc050c83",
   728 => x"ffe08c08",
   729 => x"fc050880",
   730 => x"2ebf3880",
   731 => x"5284d480",
   732 => x"c051f5bd",
   733 => x"3f83ffe0",
   734 => x"80085372",
   735 => x"812e0981",
   736 => x"068b3881",
   737 => x"0b83ffe0",
   738 => x"8c08fc05",
   739 => x"0c83ffe0",
   740 => x"8c08fc05",
   741 => x"08822e09",
   742 => x"8106ffb1",
   743 => x"38800b83",
   744 => x"ffe08c08",
   745 => x"f4050cbb",
   746 => x"39fafe3f",
   747 => x"83ffe080",
   748 => x"087083ff",
   749 => x"e1ac0c53",
   750 => x"815287fc",
   751 => x"80d051f4",
   752 => x"f03f81ff",
   753 => x"0b86e980",
   754 => x"8023830b",
   755 => x"86e98084",
   756 => x"2381ff0b",
   757 => x"86e98080",
   758 => x"23810b83",
   759 => x"ffe08c08",
   760 => x"f4050c83",
   761 => x"ffe08c08",
   762 => x"f4050883",
   763 => x"ffe0800c",
   764 => x"873d0d83",
   765 => x"ffe08c0c",
   766 => x"0483ffe0",
   767 => x"8c080283",
   768 => x"ffe08c0c",
   769 => x"803d0d80",
   770 => x"7083ffe0",
   771 => x"800c5182",
   772 => x"3d0d83ff",
   773 => x"e08c0c04",
   774 => x"83ffe08c",
   775 => x"080283ff",
   776 => x"e08c0cf5",
   777 => x"3d0d800b",
   778 => x"83ffe08c",
   779 => x"08fc050c",
   780 => x"81ff0b86",
   781 => x"e9808023",
   782 => x"820b86e9",
   783 => x"80842381",
   784 => x"0b86e980",
   785 => x"882381ff",
   786 => x"0b86e980",
   787 => x"802383ff",
   788 => x"e08c0888",
   789 => x"05085287",
   790 => x"fc80d151",
   791 => x"f3d33f83",
   792 => x"ffe08008",
   793 => x"7083ffe0",
   794 => x"8c08f405",
   795 => x"0c5483ff",
   796 => x"e08c08f4",
   797 => x"0508802e",
   798 => x"b13883ff",
   799 => x"e08c08f4",
   800 => x"05085383",
   801 => x"ffe08c08",
   802 => x"88050852",
   803 => x"848080ad",
   804 => x"d451e7f0",
   805 => x"3f83ffe0",
   806 => x"8c08fc05",
   807 => x"087083ff",
   808 => x"e08c08e0",
   809 => x"050c5481",
   810 => x"fa3980db",
   811 => x"c6e00b83",
   812 => x"ffe08c08",
   813 => x"f8050c83",
   814 => x"ffe08c08",
   815 => x"f80508ff",
   816 => x"0583ffe0",
   817 => x"8c08f805",
   818 => x"0c83ffe0",
   819 => x"8c08f805",
   820 => x"08802e81",
   821 => x"ad3881ff",
   822 => x"0b86e980",
   823 => x"802386e9",
   824 => x"80802270",
   825 => x"83ffff06",
   826 => x"7081ff06",
   827 => x"83ffe08c",
   828 => x"08f0050c",
   829 => x"515483ff",
   830 => x"e08c08f0",
   831 => x"050881fe",
   832 => x"2e098106",
   833 => x"ffb13880",
   834 => x"0b83ffe0",
   835 => x"8c08ec05",
   836 => x"0c83ffe0",
   837 => x"8c08ec05",
   838 => x"0880ff24",
   839 => x"80cd38f0",
   840 => x"b33f83ff",
   841 => x"e0800870",
   842 => x"83ffe08c",
   843 => x"08e8050c",
   844 => x"83ffe08c",
   845 => x"088c0508",
   846 => x"83ffe08c",
   847 => x"08e80508",
   848 => x"710c83ff",
   849 => x"e08c088c",
   850 => x"05088405",
   851 => x"83ffe08c",
   852 => x"088c050c",
   853 => x"83ffe08c",
   854 => x"08ec0508",
   855 => x"810583ff",
   856 => x"e08c08ec",
   857 => x"050c5154",
   858 => x"ffa73981",
   859 => x"0b83ffe0",
   860 => x"8c08f805",
   861 => x"0c810b83",
   862 => x"ffe08c08",
   863 => x"fc050cfe",
   864 => x"b63981ff",
   865 => x"0b86e980",
   866 => x"8023830b",
   867 => x"86e98084",
   868 => x"2383ffe0",
   869 => x"8c08fc05",
   870 => x"087083ff",
   871 => x"e08c08e0",
   872 => x"050c5483",
   873 => x"ffe08c08",
   874 => x"e0050883",
   875 => x"ffe0800c",
   876 => x"8d3d0d83",
   877 => x"ffe08c0c",
   878 => x"0402fc05",
   879 => x"0d7083ff",
   880 => x"e0800c02",
   881 => x"84050d04",
   882 => x"02f8050d",
   883 => x"848080ad",
   884 => x"f4518480",
   885 => x"8086dc2d",
   886 => x"84808096",
   887 => x"962d83ff",
   888 => x"e0800880",
   889 => x"2ebc3884",
   890 => x"8080ae8c",
   891 => x"51848080",
   892 => x"86dc2d84",
   893 => x"80809d86",
   894 => x"2d805284",
   895 => x"8080aea4",
   896 => x"51848080",
   897 => x"a9e92d83",
   898 => x"ffe08008",
   899 => x"802e8738",
   900 => x"84808080",
   901 => x"8c2d8480",
   902 => x"80aeb051",
   903 => x"84808086",
   904 => x"dc2d8480",
   905 => x"80aec851",
   906 => x"84808086",
   907 => x"dc2d800b",
   908 => x"83ffe080",
   909 => x"0c028805",
   910 => x"0d0402e8",
   911 => x"050d7779",
   912 => x"7b585555",
   913 => x"80537276",
   914 => x"25af3874",
   915 => x"70810556",
   916 => x"84808080",
   917 => x"af2d7470",
   918 => x"81055684",
   919 => x"808080af",
   920 => x"2d525271",
   921 => x"712e8938",
   922 => x"81518480",
   923 => x"809cfb04",
   924 => x"81135384",
   925 => x"80809cc6",
   926 => x"04805170",
   927 => x"83ffe080",
   928 => x"0c029805",
   929 => x"0d0402d8",
   930 => x"050dff0b",
   931 => x"83ffe5d8",
   932 => x"0c800b83",
   933 => x"ffe5ec0c",
   934 => x"848080ae",
   935 => x"e8518480",
   936 => x"8086dc2d",
   937 => x"83ffe1c4",
   938 => x"52805184",
   939 => x"80809898",
   940 => x"2d83ffe0",
   941 => x"80085483",
   942 => x"ffe08008",
   943 => x"95388480",
   944 => x"80aef851",
   945 => x"84808086",
   946 => x"dc2d7355",
   947 => x"848080a5",
   948 => x"ab048480",
   949 => x"80af8c51",
   950 => x"84808086",
   951 => x"dc2d8056",
   952 => x"810b83ff",
   953 => x"e1b80c88",
   954 => x"53848080",
   955 => x"afa45283",
   956 => x"ffe1fa51",
   957 => x"8480809c",
   958 => x"ba2d83ff",
   959 => x"e0800876",
   960 => x"2e098106",
   961 => x"8b3883ff",
   962 => x"e0800883",
   963 => x"ffe1b80c",
   964 => x"88538480",
   965 => x"80afb052",
   966 => x"83ffe296",
   967 => x"51848080",
   968 => x"9cba2d83",
   969 => x"ffe08008",
   970 => x"8b3883ff",
   971 => x"e0800883",
   972 => x"ffe1b80c",
   973 => x"83ffe1b8",
   974 => x"08528480",
   975 => x"80afbc51",
   976 => x"84808081",
   977 => x"842d83ff",
   978 => x"e1b80880",
   979 => x"2e81cb38",
   980 => x"83ffe58a",
   981 => x"0b848080",
   982 => x"80af2d83",
   983 => x"ffe58b0b",
   984 => x"84808080",
   985 => x"af2d7198",
   986 => x"2b71902b",
   987 => x"0783ffe5",
   988 => x"8c0b8480",
   989 => x"8080af2d",
   990 => x"70882b72",
   991 => x"0783ffe5",
   992 => x"8d0b8480",
   993 => x"8080af2d",
   994 => x"710783ff",
   995 => x"e5c20b84",
   996 => x"808080af",
   997 => x"2d83ffe5",
   998 => x"c30b8480",
   999 => x"8080af2d",
  1000 => x"71882b07",
  1001 => x"535f5452",
  1002 => x"5a565755",
  1003 => x"7381abaa",
  1004 => x"2e098106",
  1005 => x"95387551",
  1006 => x"84808083",
  1007 => x"ee2d83ff",
  1008 => x"e0800856",
  1009 => x"8480809f",
  1010 => x"e3047382",
  1011 => x"d4d52e93",
  1012 => x"38848080",
  1013 => x"afd05184",
  1014 => x"808086dc",
  1015 => x"2d848080",
  1016 => x"a1ef0475",
  1017 => x"52848080",
  1018 => x"aff05184",
  1019 => x"80808184",
  1020 => x"2d83ffe1",
  1021 => x"c4527551",
  1022 => x"84808098",
  1023 => x"982d83ff",
  1024 => x"e0800855",
  1025 => x"83ffe080",
  1026 => x"08802e85",
  1027 => x"9e388480",
  1028 => x"80b08851",
  1029 => x"84808086",
  1030 => x"dc2d8480",
  1031 => x"80b0b051",
  1032 => x"84808081",
  1033 => x"842d8853",
  1034 => x"848080af",
  1035 => x"b05283ff",
  1036 => x"e2965184",
  1037 => x"80809cba",
  1038 => x"2d83ffe0",
  1039 => x"80088e38",
  1040 => x"810b83ff",
  1041 => x"e5ec0c84",
  1042 => x"8080a0fb",
  1043 => x"04885384",
  1044 => x"8080afa4",
  1045 => x"5283ffe1",
  1046 => x"fa518480",
  1047 => x"809cba2d",
  1048 => x"83ffe080",
  1049 => x"08802e93",
  1050 => x"38848080",
  1051 => x"b0c85184",
  1052 => x"80808184",
  1053 => x"2d848080",
  1054 => x"a1ef0483",
  1055 => x"ffe5c20b",
  1056 => x"84808080",
  1057 => x"af2d5473",
  1058 => x"80d52e09",
  1059 => x"810680df",
  1060 => x"3883ffe5",
  1061 => x"c30b8480",
  1062 => x"8080af2d",
  1063 => x"547381aa",
  1064 => x"2e098106",
  1065 => x"80c93880",
  1066 => x"0b83ffe1",
  1067 => x"c40b8480",
  1068 => x"8080af2d",
  1069 => x"56547481",
  1070 => x"e92e8338",
  1071 => x"81547481",
  1072 => x"eb2e8c38",
  1073 => x"80557375",
  1074 => x"2e098106",
  1075 => x"83dd3883",
  1076 => x"ffe1cf0b",
  1077 => x"84808080",
  1078 => x"af2d5574",
  1079 => x"923883ff",
  1080 => x"e1d00b84",
  1081 => x"808080af",
  1082 => x"2d547382",
  1083 => x"2e893880",
  1084 => x"55848080",
  1085 => x"a5ab0483",
  1086 => x"ffe1d10b",
  1087 => x"84808080",
  1088 => x"af2d7083",
  1089 => x"ffe5f40c",
  1090 => x"ff0583ff",
  1091 => x"e5e80c83",
  1092 => x"ffe1d20b",
  1093 => x"84808080",
  1094 => x"af2d83ff",
  1095 => x"e1d30b84",
  1096 => x"808080af",
  1097 => x"2d587605",
  1098 => x"77828029",
  1099 => x"057083ff",
  1100 => x"e5dc0c83",
  1101 => x"ffe1d40b",
  1102 => x"84808080",
  1103 => x"af2d7083",
  1104 => x"ffe5d40c",
  1105 => x"83ffe5ec",
  1106 => x"08595758",
  1107 => x"76802e81",
  1108 => x"ea388853",
  1109 => x"848080af",
  1110 => x"b05283ff",
  1111 => x"e2965184",
  1112 => x"80809cba",
  1113 => x"2d83ffe0",
  1114 => x"800882bf",
  1115 => x"3883ffe5",
  1116 => x"f4087084",
  1117 => x"2b83ffe5",
  1118 => x"c40c7083",
  1119 => x"ffe5f00c",
  1120 => x"83ffe1e9",
  1121 => x"0b848080",
  1122 => x"80af2d83",
  1123 => x"ffe1e80b",
  1124 => x"84808080",
  1125 => x"af2d7182",
  1126 => x"80290583",
  1127 => x"ffe1ea0b",
  1128 => x"84808080",
  1129 => x"af2d7084",
  1130 => x"80802912",
  1131 => x"83ffe1eb",
  1132 => x"0b848080",
  1133 => x"80af2d70",
  1134 => x"81800a29",
  1135 => x"127083ff",
  1136 => x"e1bc0c83",
  1137 => x"ffe5d408",
  1138 => x"712983ff",
  1139 => x"e5dc0805",
  1140 => x"7083ffe5",
  1141 => x"fc0c83ff",
  1142 => x"e1f10b84",
  1143 => x"808080af",
  1144 => x"2d83ffe1",
  1145 => x"f00b8480",
  1146 => x"8080af2d",
  1147 => x"71828029",
  1148 => x"0583ffe1",
  1149 => x"f20b8480",
  1150 => x"8080af2d",
  1151 => x"70848080",
  1152 => x"291283ff",
  1153 => x"e1f30b84",
  1154 => x"808080af",
  1155 => x"2d70982b",
  1156 => x"81f00a06",
  1157 => x"72057083",
  1158 => x"ffe1c00c",
  1159 => x"fe117e29",
  1160 => x"770583ff",
  1161 => x"e5e40c52",
  1162 => x"59524354",
  1163 => x"5e515259",
  1164 => x"525d5759",
  1165 => x"57848080",
  1166 => x"a5a90483",
  1167 => x"ffe1d60b",
  1168 => x"84808080",
  1169 => x"af2d83ff",
  1170 => x"e1d50b84",
  1171 => x"808080af",
  1172 => x"2d718280",
  1173 => x"29057083",
  1174 => x"ffe5c40c",
  1175 => x"70a02983",
  1176 => x"ff057089",
  1177 => x"2a7083ff",
  1178 => x"e5f00c83",
  1179 => x"ffe1db0b",
  1180 => x"84808080",
  1181 => x"af2d83ff",
  1182 => x"e1da0b84",
  1183 => x"808080af",
  1184 => x"2d718280",
  1185 => x"29057083",
  1186 => x"ffe1bc0c",
  1187 => x"7b71291e",
  1188 => x"7083ffe5",
  1189 => x"e40c7d83",
  1190 => x"ffe1c00c",
  1191 => x"730583ff",
  1192 => x"e5fc0c55",
  1193 => x"5e515155",
  1194 => x"55815574",
  1195 => x"83ffe080",
  1196 => x"0c02a805",
  1197 => x"0d0402ec",
  1198 => x"050d7670",
  1199 => x"872c7180",
  1200 => x"ff065755",
  1201 => x"5383ffe5",
  1202 => x"ec088a38",
  1203 => x"72882c73",
  1204 => x"81ff0656",
  1205 => x"547383ff",
  1206 => x"e5d8082e",
  1207 => x"a93883ff",
  1208 => x"e1c45283",
  1209 => x"ffe5dc08",
  1210 => x"14518480",
  1211 => x"8098982d",
  1212 => x"83ffe080",
  1213 => x"085383ff",
  1214 => x"e0800880",
  1215 => x"2e80cf38",
  1216 => x"7383ffe5",
  1217 => x"d80c83ff",
  1218 => x"e5ec0880",
  1219 => x"2ea23874",
  1220 => x"842983ff",
  1221 => x"e1c40570",
  1222 => x"08525384",
  1223 => x"808083ee",
  1224 => x"2d83ffe0",
  1225 => x"8008f00a",
  1226 => x"06558480",
  1227 => x"80a6cc04",
  1228 => x"741083ff",
  1229 => x"e1c40570",
  1230 => x"84808080",
  1231 => x"9a2d5253",
  1232 => x"84808084",
  1233 => x"a02d83ff",
  1234 => x"e0800855",
  1235 => x"74537283",
  1236 => x"ffe0800c",
  1237 => x"0294050d",
  1238 => x"0402cc05",
  1239 => x"0d7e605e",
  1240 => x"5b8056ff",
  1241 => x"0b83ffe5",
  1242 => x"d80c83ff",
  1243 => x"e1c00883",
  1244 => x"ffe5e408",
  1245 => x"565783ff",
  1246 => x"e5ec0876",
  1247 => x"2e8f3883",
  1248 => x"ffe5f408",
  1249 => x"842b5984",
  1250 => x"8080a795",
  1251 => x"0483ffe5",
  1252 => x"f008842b",
  1253 => x"59805a79",
  1254 => x"792781f0",
  1255 => x"38798f06",
  1256 => x"a0175754",
  1257 => x"73a43874",
  1258 => x"52848080",
  1259 => x"b0e85184",
  1260 => x"80808184",
  1261 => x"2d83ffe1",
  1262 => x"c4527451",
  1263 => x"81155584",
  1264 => x"80809898",
  1265 => x"2d83ffe1",
  1266 => x"c4568076",
  1267 => x"84808080",
  1268 => x"af2d5558",
  1269 => x"73782e83",
  1270 => x"38815873",
  1271 => x"81e52e81",
  1272 => x"a2388170",
  1273 => x"7906555c",
  1274 => x"73802e81",
  1275 => x"96388b16",
  1276 => x"84808080",
  1277 => x"af2d9806",
  1278 => x"58778187",
  1279 => x"388b537c",
  1280 => x"52755184",
  1281 => x"80809cba",
  1282 => x"2d83ffe0",
  1283 => x"800880f3",
  1284 => x"389c1608",
  1285 => x"51848080",
  1286 => x"83ee2d83",
  1287 => x"ffe08008",
  1288 => x"841c0c9a",
  1289 => x"16848080",
  1290 => x"809a2d51",
  1291 => x"84808084",
  1292 => x"a02d83ff",
  1293 => x"e0800883",
  1294 => x"ffe08008",
  1295 => x"555583ff",
  1296 => x"e5ec0880",
  1297 => x"2ea03894",
  1298 => x"16848080",
  1299 => x"809a2d51",
  1300 => x"84808084",
  1301 => x"a02d83ff",
  1302 => x"e0800890",
  1303 => x"2b83fff0",
  1304 => x"0a067016",
  1305 => x"51547388",
  1306 => x"1c0c777b",
  1307 => x"0c7c5284",
  1308 => x"8080b188",
  1309 => x"51848080",
  1310 => x"81842d7b",
  1311 => x"54848080",
  1312 => x"a9de0481",
  1313 => x"1a5a8480",
  1314 => x"80a79704",
  1315 => x"83ffe5ec",
  1316 => x"08802e80",
  1317 => x"c7387651",
  1318 => x"848080a5",
  1319 => x"b62d83ff",
  1320 => x"e0800883",
  1321 => x"ffe08008",
  1322 => x"53848080",
  1323 => x"b19c5257",
  1324 => x"84808081",
  1325 => x"842d7680",
  1326 => x"fffffff8",
  1327 => x"06547380",
  1328 => x"fffffff8",
  1329 => x"2e9638fe",
  1330 => x"1783ffe5",
  1331 => x"f4082983",
  1332 => x"ffe5fc08",
  1333 => x"05558480",
  1334 => x"80a79504",
  1335 => x"80547383",
  1336 => x"ffe0800c",
  1337 => x"02b4050d",
  1338 => x"0402e405",
  1339 => x"0d787a71",
  1340 => x"5483ffe5",
  1341 => x"c8535555",
  1342 => x"848080a6",
  1343 => x"d92d83ff",
  1344 => x"e0800881",
  1345 => x"ff065372",
  1346 => x"802e8188",
  1347 => x"38848080",
  1348 => x"b1b45184",
  1349 => x"808086dc",
  1350 => x"2d83ffe5",
  1351 => x"cc0883ff",
  1352 => x"05892a57",
  1353 => x"80705656",
  1354 => x"75772581",
  1355 => x"873883ff",
  1356 => x"e5d008fe",
  1357 => x"0583ffe5",
  1358 => x"f4082983",
  1359 => x"ffe5fc08",
  1360 => x"117683ff",
  1361 => x"e5e80806",
  1362 => x"05755452",
  1363 => x"53848080",
  1364 => x"98982d83",
  1365 => x"ffe08008",
  1366 => x"802e80cc",
  1367 => x"38811570",
  1368 => x"83ffe5e8",
  1369 => x"08065455",
  1370 => x"72973883",
  1371 => x"ffe5d008",
  1372 => x"51848080",
  1373 => x"a5b62d83",
  1374 => x"ffe08008",
  1375 => x"83ffe5d0",
  1376 => x"0c848014",
  1377 => x"81175754",
  1378 => x"767624ff",
  1379 => x"a1388480",
  1380 => x"80abb404",
  1381 => x"74528480",
  1382 => x"80b1d051",
  1383 => x"84808081",
  1384 => x"842d8480",
  1385 => x"80abb604",
  1386 => x"83ffe080",
  1387 => x"08538480",
  1388 => x"80abb604",
  1389 => x"81537283",
  1390 => x"ffe0800c",
  1391 => x"029c050d",
  1392 => x"0483ffe0",
  1393 => x"8c080283",
  1394 => x"ffe08c0c",
  1395 => x"ff3d0d80",
  1396 => x"0b83ffe0",
  1397 => x"8c08fc05",
  1398 => x"0c83ffe0",
  1399 => x"8c088805",
  1400 => x"088106ff",
  1401 => x"11700970",
  1402 => x"83ffe08c",
  1403 => x"088c0508",
  1404 => x"0683ffe0",
  1405 => x"8c08fc05",
  1406 => x"081183ff",
  1407 => x"e08c08fc",
  1408 => x"050c83ff",
  1409 => x"e08c0888",
  1410 => x"0508812a",
  1411 => x"83ffe08c",
  1412 => x"0888050c",
  1413 => x"83ffe08c",
  1414 => x"088c0508",
  1415 => x"1083ffe0",
  1416 => x"8c088c05",
  1417 => x"0c515151",
  1418 => x"5183ffe0",
  1419 => x"8c088805",
  1420 => x"08802e84",
  1421 => x"38ffa239",
  1422 => x"83ffe08c",
  1423 => x"08fc0508",
  1424 => x"7083ffe0",
  1425 => x"800c5183",
  1426 => x"3d0d83ff",
  1427 => x"e08c0c04",
  1428 => x"00ffffff",
  1429 => x"ff00ffff",
  1430 => x"ffff00ff",
  1431 => x"ffffff00",
  1432 => x"436d645f",
  1433 => x"696e6974",
  1434 => x"0a000000",
  1435 => x"636d645f",
  1436 => x"434d4438",
  1437 => x"20726573",
  1438 => x"706f6e73",
  1439 => x"653a2025",
  1440 => x"640a0000",
  1441 => x"434d4438",
  1442 => x"5f342072",
  1443 => x"6573706f",
  1444 => x"6e73653a",
  1445 => x"2025640a",
  1446 => x"00000000",
  1447 => x"434d4435",
  1448 => x"38202564",
  1449 => x"0a202000",
  1450 => x"434d4435",
  1451 => x"385f3220",
  1452 => x"25640a20",
  1453 => x"20000000",
  1454 => x"53444843",
  1455 => x"20496e69",
  1456 => x"7469616c",
  1457 => x"697a6174",
  1458 => x"696f6e20",
  1459 => x"6572726f",
  1460 => x"72210a00",
  1461 => x"52656164",
  1462 => x"20636f6d",
  1463 => x"6d616e64",
  1464 => x"20666169",
  1465 => x"6c656420",
  1466 => x"61742025",
  1467 => x"64202825",
  1468 => x"64290a00",
  1469 => x"496e6974",
  1470 => x"69616c69",
  1471 => x"7a696e67",
  1472 => x"20534420",
  1473 => x"63617264",
  1474 => x"0a000000",
  1475 => x"48756e74",
  1476 => x"696e6720",
  1477 => x"666f7220",
  1478 => x"70617274",
  1479 => x"6974696f",
  1480 => x"6e0a0000",
  1481 => x"4f53445a",
  1482 => x"50553031",
  1483 => x"53595300",
  1484 => x"43616e27",
  1485 => x"74206c6f",
  1486 => x"61642066",
  1487 => x"69726d77",
  1488 => x"6172650a",
  1489 => x"00000000",
  1490 => x"4661696c",
  1491 => x"65642074",
  1492 => x"6f20696e",
  1493 => x"69746961",
  1494 => x"6c697a65",
  1495 => x"20534420",
  1496 => x"63617264",
  1497 => x"0a000000",
  1498 => x"52656164",
  1499 => x"696e6720",
  1500 => x"4d42520a",
  1501 => x"00000000",
  1502 => x"52656164",
  1503 => x"206f6620",
  1504 => x"4d425220",
  1505 => x"6661696c",
  1506 => x"65640a00",
  1507 => x"4d425220",
  1508 => x"73756363",
  1509 => x"65737366",
  1510 => x"756c6c79",
  1511 => x"20726561",
  1512 => x"640a0000",
  1513 => x"46415431",
  1514 => x"36202020",
  1515 => x"00000000",
  1516 => x"46415433",
  1517 => x"32202020",
  1518 => x"00000000",
  1519 => x"50617274",
  1520 => x"6974696f",
  1521 => x"6e636f75",
  1522 => x"6e742025",
  1523 => x"640a0000",
  1524 => x"4e6f2070",
  1525 => x"61727469",
  1526 => x"74696f6e",
  1527 => x"20736967",
  1528 => x"6e617475",
  1529 => x"72652066",
  1530 => x"6f756e64",
  1531 => x"0a000000",
  1532 => x"52656164",
  1533 => x"696e6720",
  1534 => x"626f6f74",
  1535 => x"20736563",
  1536 => x"746f7220",
  1537 => x"25640a00",
  1538 => x"52656164",
  1539 => x"20626f6f",
  1540 => x"74207365",
  1541 => x"63746f72",
  1542 => x"2066726f",
  1543 => x"6d206669",
  1544 => x"72737420",
  1545 => x"70617274",
  1546 => x"6974696f",
  1547 => x"6e0a0000",
  1548 => x"48756e74",
  1549 => x"696e6720",
  1550 => x"666f7220",
  1551 => x"66696c65",
  1552 => x"73797374",
  1553 => x"656d0a00",
  1554 => x"556e7375",
  1555 => x"70706f72",
  1556 => x"74656420",
  1557 => x"70617274",
  1558 => x"6974696f",
  1559 => x"6e207479",
  1560 => x"7065210d",
  1561 => x"00000000",
  1562 => x"52656164",
  1563 => x"696e6720",
  1564 => x"64697265",
  1565 => x"63746f72",
  1566 => x"79207365",
  1567 => x"63746f72",
  1568 => x"2025640a",
  1569 => x"00000000",
  1570 => x"66696c65",
  1571 => x"20222573",
  1572 => x"2220666f",
  1573 => x"756e640d",
  1574 => x"00000000",
  1575 => x"47657446",
  1576 => x"41544c69",
  1577 => x"6e6b2072",
  1578 => x"65747572",
  1579 => x"6e656420",
  1580 => x"25640a00",
  1581 => x"4f70656e",
  1582 => x"65642066",
  1583 => x"696c652c",
  1584 => x"206c6f61",
  1585 => x"64696e67",
  1586 => x"2e2e2e0a",
  1587 => x"00000000",
  1588 => x"43616e27",
  1589 => x"74206f70",
  1590 => x"656e2025",
  1591 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

