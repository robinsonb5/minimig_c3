-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity DiagROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end DiagROM_ROM;

architecture arch of DiagROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808088",
     1 => x"e8040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90088480",
    10 => x"8088e408",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b848080",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"84808088",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"09810584",
    90 => x"8080889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"84808096",
   162 => x"90738306",
   163 => x"10100508",
   164 => x"06848080",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"8480808f",
   171 => x"c62d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"84808091",
   179 => x"ee2d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"80048480",
   279 => x"8088da04",
   280 => x"04000000",
   281 => x"40000460",
   282 => x"84808088",
   283 => x"da0b8480",
   284 => x"8088f404",
   285 => x"02fc050d",
   286 => x"84808096",
   287 => x"a0518480",
   288 => x"80898a2d",
   289 => x"84808089",
   290 => x"840402d8",
   291 => x"050d7b59",
   292 => x"78802e90",
   293 => x"38788480",
   294 => x"8096b00c",
   295 => x"800b8480",
   296 => x"8096b80c",
   297 => x"84808096",
   298 => x"b8085271",
   299 => x"83813884",
   300 => x"808096b0",
   301 => x"08841184",
   302 => x"808096b0",
   303 => x"0c700884",
   304 => x"808096b4",
   305 => x"0c518112",
   306 => x"83068480",
   307 => x"8096b408",
   308 => x"70982c53",
   309 => x"5856800b",
   310 => x"84808096",
   311 => x"b0085353",
   312 => x"70802eaf",
   313 => x"38758480",
   314 => x"8096b80c",
   315 => x"81135375",
   316 => x"829e3871",
   317 => x"84137108",
   318 => x"84808096",
   319 => x"b40c8118",
   320 => x"83068480",
   321 => x"8096b408",
   322 => x"70982c55",
   323 => x"5a585354",
   324 => x"70d33871",
   325 => x"84808096",
   326 => x"b00c810b",
   327 => x"82147072",
   328 => x"2a5c5955",
   329 => x"900b86e9",
   330 => x"80842390",
   331 => x"0b86e980",
   332 => x"803486e9",
   333 => x"80803352",
   334 => x"810b86e9",
   335 => x"80803486",
   336 => x"e9808033",
   337 => x"51800b86",
   338 => x"e9808034",
   339 => x"86e98080",
   340 => x"3351800b",
   341 => x"86e98080",
   342 => x"3486e980",
   343 => x"80335180",
   344 => x"0b86e980",
   345 => x"803486e9",
   346 => x"80803370",
   347 => x"81ff0655",
   348 => x"53800b86",
   349 => x"e9808034",
   350 => x"86e98080",
   351 => x"337081ff",
   352 => x"06738106",
   353 => x"54545171",
   354 => x"802e80f7",
   355 => x"3874802e",
   356 => x"81e63873",
   357 => x"81803270",
   358 => x"09810570",
   359 => x"80255356",
   360 => x"5272862e",
   361 => x"09810681",
   362 => x"b4388170",
   363 => x"72065552",
   364 => x"73802e81",
   365 => x"a8388055",
   366 => x"fed5ca0b",
   367 => x"86e98080",
   368 => x"2386e980",
   369 => x"80225171",
   370 => x"86e98080",
   371 => x"2386e980",
   372 => x"80225174",
   373 => x"86e98080",
   374 => x"2386e980",
   375 => x"80225177",
   376 => x"86e98080",
   377 => x"2386e980",
   378 => x"80225174",
   379 => x"86e98080",
   380 => x"2386e980",
   381 => x"80225174",
   382 => x"86e98080",
   383 => x"2386e980",
   384 => x"80225191",
   385 => x"0b86e980",
   386 => x"84238480",
   387 => x"808aa404",
   388 => x"76882b84",
   389 => x"808096b4",
   390 => x"0c811683",
   391 => x"06848080",
   392 => x"96b40870",
   393 => x"982c5358",
   394 => x"56848080",
   395 => x"8a900484",
   396 => x"808096b4",
   397 => x"08882b84",
   398 => x"808096b4",
   399 => x"0c811283",
   400 => x"06848080",
   401 => x"96b40870",
   402 => x"982c5358",
   403 => x"56800b84",
   404 => x"808096b0",
   405 => x"08535384",
   406 => x"808089e0",
   407 => x"04758480",
   408 => x"8096b80c",
   409 => x"910b86e9",
   410 => x"80842380",
   411 => x"0b848080",
   412 => x"80880c02",
   413 => x"a8050d04",
   414 => x"7381802e",
   415 => x"098106dd",
   416 => x"3879732e",
   417 => x"098106d5",
   418 => x"38721053",
   419 => x"78802e81",
   420 => x"ee387884",
   421 => x"808096b0",
   422 => x"0c748480",
   423 => x"8096b80c",
   424 => x"84808096",
   425 => x"b8085271",
   426 => x"81c63884",
   427 => x"808096b0",
   428 => x"08841184",
   429 => x"808096b0",
   430 => x"0c700884",
   431 => x"808096b4",
   432 => x"0c568112",
   433 => x"83068480",
   434 => x"8096b80c",
   435 => x"84808096",
   436 => x"b4087098",
   437 => x"2cff1555",
   438 => x"535472ff",
   439 => x"2e80d938",
   440 => x"84808096",
   441 => x"b0085571",
   442 => x"86e98080",
   443 => x"3486e980",
   444 => x"80335171",
   445 => x"802eae38",
   446 => x"84808096",
   447 => x"b8085271",
   448 => x"80ca3874",
   449 => x"84167108",
   450 => x"84808096",
   451 => x"b40c8114",
   452 => x"83068480",
   453 => x"8096b80c",
   454 => x"84808096",
   455 => x"b4087098",
   456 => x"2c555656",
   457 => x"57ff1353",
   458 => x"72ff2e09",
   459 => x"8106ffb7",
   460 => x"38748480",
   461 => x"8096b00c",
   462 => x"910b86e9",
   463 => x"80842381",
   464 => x"0b848080",
   465 => x"80880c02",
   466 => x"a8050d04",
   467 => x"73882b84",
   468 => x"808096b4",
   469 => x"0c811283",
   470 => x"06848080",
   471 => x"96b80c84",
   472 => x"808096b4",
   473 => x"0870982c",
   474 => x"53548480",
   475 => x"808ea504",
   476 => x"76882b84",
   477 => x"808096b4",
   478 => x"0c848080",
   479 => x"8dc20475",
   480 => x"84808096",
   481 => x"b80c8480",
   482 => x"808da004",
   483 => x"02f0050d",
   484 => x"86e98084",
   485 => x"53907323",
   486 => x"86e98080",
   487 => x"51807123",
   488 => x"70227083",
   489 => x"ffff0653",
   490 => x"54807123",
   491 => x"70225480",
   492 => x"71237022",
   493 => x"51917323",
   494 => x"71882a84",
   495 => x"80808088",
   496 => x"0c029005",
   497 => x"0d048480",
   498 => x"80809408",
   499 => x"02848080",
   500 => x"80940cf9",
   501 => x"3d0d800b",
   502 => x"84808080",
   503 => x"9408fc05",
   504 => x"0c848080",
   505 => x"80940888",
   506 => x"05088025",
   507 => x"80c73884",
   508 => x"80808094",
   509 => x"08880508",
   510 => x"30848080",
   511 => x"80940888",
   512 => x"050c800b",
   513 => x"84808080",
   514 => x"9408f405",
   515 => x"0c848080",
   516 => x"809408fc",
   517 => x"05088c38",
   518 => x"810b8480",
   519 => x"80809408",
   520 => x"f4050c84",
   521 => x"80808094",
   522 => x"08f40508",
   523 => x"84808080",
   524 => x"9408fc05",
   525 => x"0c848080",
   526 => x"8094088c",
   527 => x"05088025",
   528 => x"80c73884",
   529 => x"80808094",
   530 => x"088c0508",
   531 => x"30848080",
   532 => x"8094088c",
   533 => x"050c800b",
   534 => x"84808080",
   535 => x"9408f005",
   536 => x"0c848080",
   537 => x"809408fc",
   538 => x"05088c38",
   539 => x"810b8480",
   540 => x"80809408",
   541 => x"f0050c84",
   542 => x"80808094",
   543 => x"08f00508",
   544 => x"84808080",
   545 => x"9408fc05",
   546 => x"0c805384",
   547 => x"80808094",
   548 => x"088c0508",
   549 => x"52848080",
   550 => x"80940888",
   551 => x"05085182",
   552 => x"983f8480",
   553 => x"80808808",
   554 => x"70848080",
   555 => x"809408f8",
   556 => x"050c5484",
   557 => x"80808094",
   558 => x"08fc0508",
   559 => x"802e9438",
   560 => x"84808080",
   561 => x"9408f805",
   562 => x"08308480",
   563 => x"80809408",
   564 => x"f8050c84",
   565 => x"80808094",
   566 => x"08f80508",
   567 => x"70848080",
   568 => x"80880c54",
   569 => x"893d0d84",
   570 => x"80808094",
   571 => x"0c048480",
   572 => x"80809408",
   573 => x"02848080",
   574 => x"80940cfb",
   575 => x"3d0d800b",
   576 => x"84808080",
   577 => x"9408fc05",
   578 => x"0c848080",
   579 => x"80940888",
   580 => x"05088025",
   581 => x"9f388480",
   582 => x"80809408",
   583 => x"88050830",
   584 => x"84808080",
   585 => x"94088805",
   586 => x"0c810b84",
   587 => x"80808094",
   588 => x"08fc050c",
   589 => x"84808080",
   590 => x"94088c05",
   591 => x"08802594",
   592 => x"38848080",
   593 => x"8094088c",
   594 => x"05083084",
   595 => x"80808094",
   596 => x"088c050c",
   597 => x"81538480",
   598 => x"80809408",
   599 => x"8c050852",
   600 => x"84808080",
   601 => x"94088805",
   602 => x"085180cd",
   603 => x"3f848080",
   604 => x"80880870",
   605 => x"84808080",
   606 => x"9408f805",
   607 => x"0c548480",
   608 => x"80809408",
   609 => x"fc050880",
   610 => x"2e943884",
   611 => x"80808094",
   612 => x"08f80508",
   613 => x"30848080",
   614 => x"809408f8",
   615 => x"050c8480",
   616 => x"80809408",
   617 => x"f8050870",
   618 => x"84808080",
   619 => x"880c5487",
   620 => x"3d0d8480",
   621 => x"8080940c",
   622 => x"04848080",
   623 => x"80940802",
   624 => x"84808080",
   625 => x"940cfd3d",
   626 => x"0d810b84",
   627 => x"80808094",
   628 => x"08fc050c",
   629 => x"800b8480",
   630 => x"80809408",
   631 => x"f8050c84",
   632 => x"80808094",
   633 => x"088c0508",
   634 => x"84808080",
   635 => x"94088805",
   636 => x"082780c5",
   637 => x"38848080",
   638 => x"809408fc",
   639 => x"0508802e",
   640 => x"b838800b",
   641 => x"84808080",
   642 => x"94088c05",
   643 => x"0824aa38",
   644 => x"84808080",
   645 => x"94088c05",
   646 => x"08108480",
   647 => x"80809408",
   648 => x"8c050c84",
   649 => x"80808094",
   650 => x"08fc0508",
   651 => x"10848080",
   652 => x"809408fc",
   653 => x"050cffa7",
   654 => x"39848080",
   655 => x"809408fc",
   656 => x"0508802e",
   657 => x"80f93884",
   658 => x"80808094",
   659 => x"088c0508",
   660 => x"84808080",
   661 => x"94088805",
   662 => x"0826b938",
   663 => x"84808080",
   664 => x"94088805",
   665 => x"08848080",
   666 => x"8094088c",
   667 => x"05083184",
   668 => x"80808094",
   669 => x"0888050c",
   670 => x"84808080",
   671 => x"9408f805",
   672 => x"08848080",
   673 => x"809408fc",
   674 => x"05080784",
   675 => x"80808094",
   676 => x"08f8050c",
   677 => x"84808080",
   678 => x"9408fc05",
   679 => x"08812a84",
   680 => x"80808094",
   681 => x"08fc050c",
   682 => x"84808080",
   683 => x"94088c05",
   684 => x"08812a84",
   685 => x"80808094",
   686 => x"088c050c",
   687 => x"fefb3984",
   688 => x"80808094",
   689 => x"08900508",
   690 => x"802e9738",
   691 => x"84808080",
   692 => x"94088805",
   693 => x"08708480",
   694 => x"80809408",
   695 => x"f4050c51",
   696 => x"95398480",
   697 => x"80809408",
   698 => x"f8050870",
   699 => x"84808080",
   700 => x"9408f405",
   701 => x"0c518480",
   702 => x"80809408",
   703 => x"f4050884",
   704 => x"80808088",
   705 => x"0c853d0d",
   706 => x"84808080",
   707 => x"940c0400",
   708 => x"00ffffff",
   709 => x"ff00ffff",
   710 => x"ffff00ff",
   711 => x"ffffff00",
   712 => x"48656c6c",
   713 => x"6f2c2077",
   714 => x"6f726c64",
   715 => x"210a0064",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

