-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity DiagROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end DiagROM_ROM;

architecture arch of DiagROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808088",
     1 => x"e8040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90088480",
    10 => x"8088e408",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b848080",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"84808088",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"09810584",
    90 => x"8080889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"84808093",
   162 => x"88738306",
   163 => x"10100508",
   164 => x"06848080",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"8480808c",
   171 => x"bc2d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"8480808e",
   179 => x"e42d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"80048480",
   279 => x"8088da04",
   280 => x"04000000",
   281 => x"40000460",
   282 => x"84808088",
   283 => x"da0b8480",
   284 => x"8088f404",
   285 => x"02fc050d",
   286 => x"84808093",
   287 => x"98518480",
   288 => x"80898a2d",
   289 => x"84808089",
   290 => x"840402e4",
   291 => x"050d7856",
   292 => x"75802e90",
   293 => x"38758480",
   294 => x"8093a80c",
   295 => x"800b8480",
   296 => x"8093b00c",
   297 => x"84808093",
   298 => x"b0085271",
   299 => x"82a93884",
   300 => x"808093a8",
   301 => x"08841184",
   302 => x"808093a8",
   303 => x"0c700884",
   304 => x"808093ac",
   305 => x"0c518112",
   306 => x"83068480",
   307 => x"8093ac08",
   308 => x"70982c84",
   309 => x"808093a8",
   310 => x"08565355",
   311 => x"5270802e",
   312 => x"ac387184",
   313 => x"808093b0",
   314 => x"0c7181cc",
   315 => x"38728414",
   316 => x"71088480",
   317 => x"8093ac0c",
   318 => x"81148306",
   319 => x"84808093",
   320 => x"ac087098",
   321 => x"2c555354",
   322 => x"545470d6",
   323 => x"38728480",
   324 => x"8093a80c",
   325 => x"900b86e9",
   326 => x"80842390",
   327 => x"0b86e980",
   328 => x"803486e9",
   329 => x"80803351",
   330 => x"810b86e9",
   331 => x"80803486",
   332 => x"e9808033",
   333 => x"51800b86",
   334 => x"e9808023",
   335 => x"86e98080",
   336 => x"2251800b",
   337 => x"86e98080",
   338 => x"3486e980",
   339 => x"80335180",
   340 => x"0b86e980",
   341 => x"803486e9",
   342 => x"80803351",
   343 => x"910b86e9",
   344 => x"80842390",
   345 => x"0b86e980",
   346 => x"8423900b",
   347 => x"86e98080",
   348 => x"3486e980",
   349 => x"80335181",
   350 => x"0b86e980",
   351 => x"803486e9",
   352 => x"80803351",
   353 => x"800b86e9",
   354 => x"80802386",
   355 => x"e9808022",
   356 => x"51800b86",
   357 => x"e9808034",
   358 => x"86e98080",
   359 => x"3351800b",
   360 => x"86e98080",
   361 => x"3486e980",
   362 => x"80335191",
   363 => x"0b86e980",
   364 => x"84238480",
   365 => x"808a9404",
   366 => x"73882b84",
   367 => x"808093ac",
   368 => x"0c811283",
   369 => x"06848080",
   370 => x"93ac0870",
   371 => x"982c5355",
   372 => x"52848080",
   373 => x"8a8a0484",
   374 => x"808093ac",
   375 => x"08882b84",
   376 => x"808093ac",
   377 => x"0c811283",
   378 => x"06848080",
   379 => x"93ac0870",
   380 => x"982c8480",
   381 => x"8093a808",
   382 => x"56535552",
   383 => x"84808089",
   384 => x"dd0402f0",
   385 => x"050d86e9",
   386 => x"80845390",
   387 => x"732386e9",
   388 => x"80805180",
   389 => x"71237022",
   390 => x"7083ffff",
   391 => x"06535480",
   392 => x"71237022",
   393 => x"54807123",
   394 => x"70225191",
   395 => x"73237188",
   396 => x"2a848080",
   397 => x"80880c02",
   398 => x"90050d04",
   399 => x"84808080",
   400 => x"94080284",
   401 => x"80808094",
   402 => x"0cf93d0d",
   403 => x"800b8480",
   404 => x"80809408",
   405 => x"fc050c84",
   406 => x"80808094",
   407 => x"08880508",
   408 => x"802580c7",
   409 => x"38848080",
   410 => x"80940888",
   411 => x"05083084",
   412 => x"80808094",
   413 => x"0888050c",
   414 => x"800b8480",
   415 => x"80809408",
   416 => x"f4050c84",
   417 => x"80808094",
   418 => x"08fc0508",
   419 => x"8c38810b",
   420 => x"84808080",
   421 => x"9408f405",
   422 => x"0c848080",
   423 => x"809408f4",
   424 => x"05088480",
   425 => x"80809408",
   426 => x"fc050c84",
   427 => x"80808094",
   428 => x"088c0508",
   429 => x"802580c7",
   430 => x"38848080",
   431 => x"8094088c",
   432 => x"05083084",
   433 => x"80808094",
   434 => x"088c050c",
   435 => x"800b8480",
   436 => x"80809408",
   437 => x"f0050c84",
   438 => x"80808094",
   439 => x"08fc0508",
   440 => x"8c38810b",
   441 => x"84808080",
   442 => x"9408f005",
   443 => x"0c848080",
   444 => x"809408f0",
   445 => x"05088480",
   446 => x"80809408",
   447 => x"fc050c80",
   448 => x"53848080",
   449 => x"8094088c",
   450 => x"05085284",
   451 => x"80808094",
   452 => x"08880508",
   453 => x"5182983f",
   454 => x"84808080",
   455 => x"88087084",
   456 => x"80808094",
   457 => x"08f8050c",
   458 => x"54848080",
   459 => x"809408fc",
   460 => x"0508802e",
   461 => x"94388480",
   462 => x"80809408",
   463 => x"f8050830",
   464 => x"84808080",
   465 => x"9408f805",
   466 => x"0c848080",
   467 => x"809408f8",
   468 => x"05087084",
   469 => x"80808088",
   470 => x"0c54893d",
   471 => x"0d848080",
   472 => x"80940c04",
   473 => x"84808080",
   474 => x"94080284",
   475 => x"80808094",
   476 => x"0cfb3d0d",
   477 => x"800b8480",
   478 => x"80809408",
   479 => x"fc050c84",
   480 => x"80808094",
   481 => x"08880508",
   482 => x"80259f38",
   483 => x"84808080",
   484 => x"94088805",
   485 => x"08308480",
   486 => x"80809408",
   487 => x"88050c81",
   488 => x"0b848080",
   489 => x"809408fc",
   490 => x"050c8480",
   491 => x"80809408",
   492 => x"8c050880",
   493 => x"25943884",
   494 => x"80808094",
   495 => x"088c0508",
   496 => x"30848080",
   497 => x"8094088c",
   498 => x"050c8153",
   499 => x"84808080",
   500 => x"94088c05",
   501 => x"08528480",
   502 => x"80809408",
   503 => x"88050851",
   504 => x"80cd3f84",
   505 => x"80808088",
   506 => x"08708480",
   507 => x"80809408",
   508 => x"f8050c54",
   509 => x"84808080",
   510 => x"9408fc05",
   511 => x"08802e94",
   512 => x"38848080",
   513 => x"809408f8",
   514 => x"05083084",
   515 => x"80808094",
   516 => x"08f8050c",
   517 => x"84808080",
   518 => x"9408f805",
   519 => x"08708480",
   520 => x"8080880c",
   521 => x"54873d0d",
   522 => x"84808080",
   523 => x"940c0484",
   524 => x"80808094",
   525 => x"08028480",
   526 => x"8080940c",
   527 => x"fd3d0d81",
   528 => x"0b848080",
   529 => x"809408fc",
   530 => x"050c800b",
   531 => x"84808080",
   532 => x"9408f805",
   533 => x"0c848080",
   534 => x"8094088c",
   535 => x"05088480",
   536 => x"80809408",
   537 => x"88050827",
   538 => x"80c53884",
   539 => x"80808094",
   540 => x"08fc0508",
   541 => x"802eb838",
   542 => x"800b8480",
   543 => x"80809408",
   544 => x"8c050824",
   545 => x"aa388480",
   546 => x"80809408",
   547 => x"8c050810",
   548 => x"84808080",
   549 => x"94088c05",
   550 => x"0c848080",
   551 => x"809408fc",
   552 => x"05081084",
   553 => x"80808094",
   554 => x"08fc050c",
   555 => x"ffa73984",
   556 => x"80808094",
   557 => x"08fc0508",
   558 => x"802e80f9",
   559 => x"38848080",
   560 => x"8094088c",
   561 => x"05088480",
   562 => x"80809408",
   563 => x"88050826",
   564 => x"b9388480",
   565 => x"80809408",
   566 => x"88050884",
   567 => x"80808094",
   568 => x"088c0508",
   569 => x"31848080",
   570 => x"80940888",
   571 => x"050c8480",
   572 => x"80809408",
   573 => x"f8050884",
   574 => x"80808094",
   575 => x"08fc0508",
   576 => x"07848080",
   577 => x"809408f8",
   578 => x"050c8480",
   579 => x"80809408",
   580 => x"fc050881",
   581 => x"2a848080",
   582 => x"809408fc",
   583 => x"050c8480",
   584 => x"80809408",
   585 => x"8c050881",
   586 => x"2a848080",
   587 => x"8094088c",
   588 => x"050cfefb",
   589 => x"39848080",
   590 => x"80940890",
   591 => x"0508802e",
   592 => x"97388480",
   593 => x"80809408",
   594 => x"88050870",
   595 => x"84808080",
   596 => x"9408f405",
   597 => x"0c519539",
   598 => x"84808080",
   599 => x"9408f805",
   600 => x"08708480",
   601 => x"80809408",
   602 => x"f4050c51",
   603 => x"84808080",
   604 => x"9408f405",
   605 => x"08848080",
   606 => x"80880c85",
   607 => x"3d0d8480",
   608 => x"8080940c",
   609 => x"04000000",
   610 => x"00ffffff",
   611 => x"ff00ffff",
   612 => x"ffff00ff",
   613 => x"ffffff00",
   614 => x"48656c6c",
   615 => x"6f2c2077",
   616 => x"6f726c64",
   617 => x"210a0064",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

