-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity DiagROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end DiagROM_ROM;

architecture arch of DiagROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ee040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"88080d80",
     5 => x"04848080",
     6 => x"80950471",
     7 => x"fd060872",
     8 => x"83060981",
     9 => x"05820583",
    10 => x"2b2a83ff",
    11 => x"ff065204",
    12 => x"71fc0608",
    13 => x"72830609",
    14 => x"81058305",
    15 => x"1010102a",
    16 => x"81ff0652",
    17 => x"0471fc06",
    18 => x"08848080",
    19 => x"9fd47383",
    20 => x"06101005",
    21 => x"08067381",
    22 => x"ff067383",
    23 => x"06098105",
    24 => x"83051010",
    25 => x"102b0772",
    26 => x"fc060c51",
    27 => x"51040284",
    28 => x"05848080",
    29 => x"80880c84",
    30 => x"80808095",
    31 => x"0b848080",
    32 => x"8fd80400",
    33 => x"02c4050d",
    34 => x"0280c005",
    35 => x"9fe0e05b",
    36 => x"56807670",
    37 => x"84055808",
    38 => x"715e5e57",
    39 => x"7c708405",
    40 => x"5e085880",
    41 => x"5b77982a",
    42 => x"78882b59",
    43 => x"54738938",
    44 => x"765e8480",
    45 => x"8083e204",
    46 => x"7b802e81",
    47 => x"fd38805c",
    48 => x"7380e42e",
    49 => x"a1387380",
    50 => x"e4268e38",
    51 => x"7380e32e",
    52 => x"819a3884",
    53 => x"808082fa",
    54 => x"047380f3",
    55 => x"2e80f538",
    56 => x"84808082",
    57 => x"fa047584",
    58 => x"1771087e",
    59 => x"5c555752",
    60 => x"7280258e",
    61 => x"38ad5184",
    62 => x"80808fca",
    63 => x"2d720981",
    64 => x"05537280",
    65 => x"2ebe3887",
    66 => x"55729c2a",
    67 => x"73842b54",
    68 => x"5271802e",
    69 => x"83388159",
    70 => x"8972258a",
    71 => x"38b71252",
    72 => x"84808082",
    73 => x"a904b012",
    74 => x"5278802e",
    75 => x"89387151",
    76 => x"8480808f",
    77 => x"ca2dff15",
    78 => x"55748025",
    79 => x"cc388480",
    80 => x"8082cc04",
    81 => x"b0518480",
    82 => x"808fca2d",
    83 => x"80538480",
    84 => x"80839304",
    85 => x"75841771",
    86 => x"0870545c",
    87 => x"57528480",
    88 => x"8085a92d",
    89 => x"7b538480",
    90 => x"80839304",
    91 => x"75841771",
    92 => x"08565752",
    93 => x"84808083",
    94 => x"ca04a551",
    95 => x"8480808f",
    96 => x"ca2d7351",
    97 => x"8480808f",
    98 => x"ca2d8217",
    99 => x"57848080",
   100 => x"83d50472",
   101 => x"ff145452",
   102 => x"807225b9",
   103 => x"38797081",
   104 => x"055b8480",
   105 => x"8080b02d",
   106 => x"70525484",
   107 => x"80808fca",
   108 => x"2d811757",
   109 => x"84808083",
   110 => x"930473a5",
   111 => x"2e098106",
   112 => x"8938815c",
   113 => x"84808083",
   114 => x"d5047351",
   115 => x"8480808f",
   116 => x"ca2d8117",
   117 => x"57811b5b",
   118 => x"837b25fd",
   119 => x"c83873fd",
   120 => x"bb387d9f",
   121 => x"e0800c02",
   122 => x"bc050d04",
   123 => x"02f4050d",
   124 => x"7470882a",
   125 => x"83fe8006",
   126 => x"7072982a",
   127 => x"0772882b",
   128 => x"87fc8080",
   129 => x"0673982b",
   130 => x"81f00a06",
   131 => x"71730707",
   132 => x"9fe0800c",
   133 => x"56515351",
   134 => x"028c050d",
   135 => x"0402f805",
   136 => x"0d028e05",
   137 => x"84808080",
   138 => x"b02d7488",
   139 => x"2b077083",
   140 => x"ffff069f",
   141 => x"e0800c51",
   142 => x"0288050d",
   143 => x"0402f805",
   144 => x"0d737090",
   145 => x"2b71902a",
   146 => x"079fe080",
   147 => x"0c520288",
   148 => x"050d0402",
   149 => x"f8050d73",
   150 => x"5170802e",
   151 => x"8c38709f",
   152 => x"e1a00c80",
   153 => x"0b9fe1a8",
   154 => x"0c9fe1a8",
   155 => x"08527198",
   156 => x"389fe1a0",
   157 => x"0884119f",
   158 => x"e1a00c70",
   159 => x"089fe1a4",
   160 => x"0c518480",
   161 => x"80859204",
   162 => x"9fe1a408",
   163 => x"882b9fe1",
   164 => x"a40c8112",
   165 => x"83069fe1",
   166 => x"a80c9fe1",
   167 => x"a408982c",
   168 => x"9fe0800c",
   169 => x"0288050d",
   170 => x"0402e805",
   171 => x"0d777052",
   172 => x"56848080",
   173 => x"84d32d9f",
   174 => x"e0800852",
   175 => x"80537180",
   176 => x"2e973881",
   177 => x"13538051",
   178 => x"84808084",
   179 => x"d32d9fe0",
   180 => x"80085284",
   181 => x"808085be",
   182 => x"04821354",
   183 => x"8155900b",
   184 => x"86e98084",
   185 => x"23a0810b",
   186 => x"86e98080",
   187 => x"2386e980",
   188 => x"80225280",
   189 => x"0b86e980",
   190 => x"802386e9",
   191 => x"80802253",
   192 => x"800b86e9",
   193 => x"80802386",
   194 => x"e9808022",
   195 => x"7083ffff",
   196 => x"0673882a",
   197 => x"70810651",
   198 => x"54515371",
   199 => x"802e81a4",
   200 => x"3874802e",
   201 => x"80e03872",
   202 => x"8280862e",
   203 => x"09810681",
   204 => x"93388055",
   205 => x"fed5ca0b",
   206 => x"86e98080",
   207 => x"2386e980",
   208 => x"80225281",
   209 => x"0b86e980",
   210 => x"802386e9",
   211 => x"80802252",
   212 => x"7486e980",
   213 => x"802386e9",
   214 => x"80802252",
   215 => x"7386e980",
   216 => x"802386e9",
   217 => x"80802252",
   218 => x"7486e980",
   219 => x"802386e9",
   220 => x"80802252",
   221 => x"7486e980",
   222 => x"802386e9",
   223 => x"80802252",
   224 => x"84808087",
   225 => x"c4047381",
   226 => x"2a828080",
   227 => x"07527272",
   228 => x"2e098106",
   229 => x"af387551",
   230 => x"84808084",
   231 => x"d32d9fe0",
   232 => x"800853ff",
   233 => x"145473ff",
   234 => x"2ea73872",
   235 => x"86e98080",
   236 => x"3486e980",
   237 => x"80335272",
   238 => x"802ee838",
   239 => x"80518480",
   240 => x"80879804",
   241 => x"910b86e9",
   242 => x"80842384",
   243 => x"808085de",
   244 => x"04910b86",
   245 => x"e9808423",
   246 => x"810b9fe0",
   247 => x"800c0298",
   248 => x"050d0402",
   249 => x"f4050d86",
   250 => x"e9808052",
   251 => x"81ff7223",
   252 => x"71225381",
   253 => x"ff722372",
   254 => x"882b83fe",
   255 => x"80067222",
   256 => x"7081ff06",
   257 => x"51525381",
   258 => x"ff722372",
   259 => x"7107882b",
   260 => x"72227081",
   261 => x"ff065152",
   262 => x"5381ff72",
   263 => x"23727107",
   264 => x"882b7222",
   265 => x"7081ff06",
   266 => x"72079fe0",
   267 => x"800c5253",
   268 => x"028c050d",
   269 => x"0402f405",
   270 => x"0d747671",
   271 => x"81ff0653",
   272 => x"53537086",
   273 => x"e9808023",
   274 => x"9fe1ac08",
   275 => x"85387189",
   276 => x"2b527198",
   277 => x"2a517086",
   278 => x"e9808023",
   279 => x"71902a70",
   280 => x"81ff0651",
   281 => x"517086e9",
   282 => x"80802371",
   283 => x"882a7081",
   284 => x"ff065151",
   285 => x"7086e980",
   286 => x"80237181",
   287 => x"ff065170",
   288 => x"86e98080",
   289 => x"2372902a",
   290 => x"7081ff06",
   291 => x"51517086",
   292 => x"e9808023",
   293 => x"86e98080",
   294 => x"227081ff",
   295 => x"06515182",
   296 => x"b8bf5270",
   297 => x"81ff2e09",
   298 => x"81069a38",
   299 => x"81ff0b86",
   300 => x"e9808023",
   301 => x"86e98080",
   302 => x"227081ff",
   303 => x"06ff1454",
   304 => x"515171df",
   305 => x"38709fe0",
   306 => x"800c028c",
   307 => x"050d0402",
   308 => x"fc050d81",
   309 => x"c75181ff",
   310 => x"0b86e980",
   311 => x"8023ff11",
   312 => x"51708025",
   313 => x"f1380284",
   314 => x"050d0402",
   315 => x"f0050d84",
   316 => x"808089cf",
   317 => x"2d819c9f",
   318 => x"53805287",
   319 => x"fc80f751",
   320 => x"84808088",
   321 => x"b52d9fe0",
   322 => x"8008549f",
   323 => x"e0800881",
   324 => x"2e098106",
   325 => x"b33881ff",
   326 => x"0b86e980",
   327 => x"8023820a",
   328 => x"52849c80",
   329 => x"e9518480",
   330 => x"8088b52d",
   331 => x"9fe08008",
   332 => x"913881ff",
   333 => x"0b86e980",
   334 => x"80237353",
   335 => x"8480808a",
   336 => x"cf048480",
   337 => x"8089cf2d",
   338 => x"ff135372",
   339 => x"ffab3872",
   340 => x"9fe0800c",
   341 => x"0290050d",
   342 => x"0402f405",
   343 => x"0d81ff0b",
   344 => x"86e98080",
   345 => x"23848080",
   346 => x"9fe45184",
   347 => x"808085a9",
   348 => x"2d935380",
   349 => x"5287fc80",
   350 => x"c1518480",
   351 => x"8088b52d",
   352 => x"9fe08008",
   353 => x"913881ff",
   354 => x"0b86e980",
   355 => x"80238153",
   356 => x"8480808b",
   357 => x"a2048480",
   358 => x"8089cf2d",
   359 => x"ff135372",
   360 => x"d238729f",
   361 => x"e0800c02",
   362 => x"8c050d04",
   363 => x"02f0050d",
   364 => x"84808089",
   365 => x"cf2d83aa",
   366 => x"52849c80",
   367 => x"c8518480",
   368 => x"8088b52d",
   369 => x"9fe08008",
   370 => x"812e0981",
   371 => x"06963884",
   372 => x"808087e3",
   373 => x"2d9fe080",
   374 => x"0883ffff",
   375 => x"06537283",
   376 => x"aa2e9d38",
   377 => x"8480808a",
   378 => x"d92d8480",
   379 => x"808bf804",
   380 => x"81548480",
   381 => x"808d8204",
   382 => x"80548480",
   383 => x"808d8204",
   384 => x"81ff0b86",
   385 => x"e9808023",
   386 => x"b1538480",
   387 => x"8089eb2d",
   388 => x"9fe08008",
   389 => x"802e80db",
   390 => x"38805287",
   391 => x"fc80fa51",
   392 => x"84808088",
   393 => x"b52d9fe0",
   394 => x"800880c7",
   395 => x"3881ff0b",
   396 => x"86e98080",
   397 => x"2386e980",
   398 => x"80225381",
   399 => x"ff0b86e9",
   400 => x"80802381",
   401 => x"ff0b86e9",
   402 => x"80802381",
   403 => x"ff0b86e9",
   404 => x"80802381",
   405 => x"ff0b86e9",
   406 => x"80802372",
   407 => x"862a7081",
   408 => x"069fe080",
   409 => x"08565153",
   410 => x"72802e96",
   411 => x"38848080",
   412 => x"8bf00472",
   413 => x"822eff80",
   414 => x"38ff1353",
   415 => x"72ff8b38",
   416 => x"7254739f",
   417 => x"e0800c02",
   418 => x"90050d04",
   419 => x"02f4050d",
   420 => x"810b9fe1",
   421 => x"ac0ca00b",
   422 => x"86e98088",
   423 => x"23830b86",
   424 => x"e9808423",
   425 => x"84808089",
   426 => x"cf2d820b",
   427 => x"86e98084",
   428 => x"23875380",
   429 => x"5284d480",
   430 => x"c0518480",
   431 => x"8088b52d",
   432 => x"9fe08008",
   433 => x"812e9738",
   434 => x"72822e09",
   435 => x"81068938",
   436 => x"80538480",
   437 => x"808e9204",
   438 => x"ff135372",
   439 => x"d6388480",
   440 => x"808bac2d",
   441 => x"9fe08008",
   442 => x"9fe1ac0c",
   443 => x"815287fc",
   444 => x"80d05184",
   445 => x"808088b5",
   446 => x"2d81ff0b",
   447 => x"86e98080",
   448 => x"23830b86",
   449 => x"e9808423",
   450 => x"81ff0b86",
   451 => x"e9808023",
   452 => x"8153729f",
   453 => x"e0800c02",
   454 => x"8c050d04",
   455 => x"800b9fe0",
   456 => x"800c0402",
   457 => x"e8050d78",
   458 => x"56805581",
   459 => x"ff0b86e9",
   460 => x"80802382",
   461 => x"0b86e980",
   462 => x"8423810b",
   463 => x"86e98088",
   464 => x"2381ff0b",
   465 => x"86e98080",
   466 => x"23775287",
   467 => x"fc80d151",
   468 => x"84808088",
   469 => x"b52d7453",
   470 => x"9fe08008",
   471 => x"752e0981",
   472 => x"0680dd38",
   473 => x"80dbc6df",
   474 => x"5481ff0b",
   475 => x"86e98080",
   476 => x"2386e980",
   477 => x"80227081",
   478 => x"ff065153",
   479 => x"7281fe2e",
   480 => x"098106a4",
   481 => x"3880ff53",
   482 => x"84808087",
   483 => x"e32d9fe0",
   484 => x"80087670",
   485 => x"8405580c",
   486 => x"ff135372",
   487 => x"8025e938",
   488 => x"81558480",
   489 => x"808faf04",
   490 => x"ff145473",
   491 => x"ffbb3881",
   492 => x"ff0b86e9",
   493 => x"80802383",
   494 => x"0b86e980",
   495 => x"84237453",
   496 => x"729fe080",
   497 => x"0c029805",
   498 => x"0d0402fc",
   499 => x"050d709f",
   500 => x"e0800c02",
   501 => x"84050d04",
   502 => x"02f8050d",
   503 => x"8480809f",
   504 => x"f0518480",
   505 => x"8085a92d",
   506 => x"8480808d",
   507 => x"8c2d9fe0",
   508 => x"8008802e",
   509 => x"bb388480",
   510 => x"80a08851",
   511 => x"84808085",
   512 => x"a92d8480",
   513 => x"8091922d",
   514 => x"80528480",
   515 => x"80a0a051",
   516 => x"8480809d",
   517 => x"892d9fe0",
   518 => x"8008802e",
   519 => x"87388480",
   520 => x"80808c2d",
   521 => x"848080a0",
   522 => x"ac518480",
   523 => x"8085a92d",
   524 => x"848080a0",
   525 => x"c4518480",
   526 => x"8085a92d",
   527 => x"800b9fe0",
   528 => x"800c0288",
   529 => x"050d0402",
   530 => x"e8050d77",
   531 => x"797b5855",
   532 => x"55805372",
   533 => x"7625af38",
   534 => x"74708105",
   535 => x"56848080",
   536 => x"80b02d74",
   537 => x"70810556",
   538 => x"84808080",
   539 => x"b02d5252",
   540 => x"71712e89",
   541 => x"38815184",
   542 => x"80809188",
   543 => x"04811353",
   544 => x"84808090",
   545 => x"d3048051",
   546 => x"709fe080",
   547 => x"0c029805",
   548 => x"0d0402d8",
   549 => x"050dff0b",
   550 => x"9fe5d80c",
   551 => x"800b9fe5",
   552 => x"ec0c8480",
   553 => x"80a0e451",
   554 => x"84808085",
   555 => x"a92d9fe1",
   556 => x"c4528051",
   557 => x"8480808e",
   558 => x"a32d9fe0",
   559 => x"8008549f",
   560 => x"e0800895",
   561 => x"38848080",
   562 => x"a0f45184",
   563 => x"808085a9",
   564 => x"2d735584",
   565 => x"808098ed",
   566 => x"04848080",
   567 => x"a1885184",
   568 => x"808085a9",
   569 => x"2d805681",
   570 => x"0b9fe1b8",
   571 => x"0c885384",
   572 => x"8080a1a0",
   573 => x"529fe1fa",
   574 => x"51848080",
   575 => x"90c72d9f",
   576 => x"e0800876",
   577 => x"2e098106",
   578 => x"89389fe0",
   579 => x"80089fe1",
   580 => x"b80c8853",
   581 => x"848080a1",
   582 => x"ac529fe2",
   583 => x"96518480",
   584 => x"8090c72d",
   585 => x"9fe08008",
   586 => x"89389fe0",
   587 => x"80089fe1",
   588 => x"b80c9fe1",
   589 => x"b8085284",
   590 => x"8080a1b8",
   591 => x"51848080",
   592 => x"81842d9f",
   593 => x"e1b80880",
   594 => x"2e81c138",
   595 => x"9fe58a0b",
   596 => x"84808080",
   597 => x"b02d9fe5",
   598 => x"8b0b8480",
   599 => x"8080b02d",
   600 => x"71982b71",
   601 => x"902b079f",
   602 => x"e58c0b84",
   603 => x"808080b0",
   604 => x"2d70882b",
   605 => x"72079fe5",
   606 => x"8d0b8480",
   607 => x"8080b02d",
   608 => x"71079fe5",
   609 => x"c20b8480",
   610 => x"8080b02d",
   611 => x"9fe5c30b",
   612 => x"84808080",
   613 => x"b02d7188",
   614 => x"2b07535f",
   615 => x"54525a56",
   616 => x"57557381",
   617 => x"abaa2e09",
   618 => x"81069438",
   619 => x"75518480",
   620 => x"8083ec2d",
   621 => x"9fe08008",
   622 => x"56848080",
   623 => x"93d80473",
   624 => x"82d4d52e",
   625 => x"93388480",
   626 => x"80a1cc51",
   627 => x"84808085",
   628 => x"a92d8480",
   629 => x"8095d704",
   630 => x"75528480",
   631 => x"80a1ec51",
   632 => x"84808081",
   633 => x"842d9fe1",
   634 => x"c4527551",
   635 => x"8480808e",
   636 => x"a32d9fe0",
   637 => x"8008559f",
   638 => x"e0800880",
   639 => x"2e84ee38",
   640 => x"848080a2",
   641 => x"84518480",
   642 => x"8085a92d",
   643 => x"848080a2",
   644 => x"ac518480",
   645 => x"8081842d",
   646 => x"88538480",
   647 => x"80a1ac52",
   648 => x"9fe29651",
   649 => x"84808090",
   650 => x"c72d9fe0",
   651 => x"80088d38",
   652 => x"810b9fe5",
   653 => x"ec0c8480",
   654 => x"8094e804",
   655 => x"88538480",
   656 => x"80a1a052",
   657 => x"9fe1fa51",
   658 => x"84808090",
   659 => x"c72d9fe0",
   660 => x"8008802e",
   661 => x"93388480",
   662 => x"80a2c451",
   663 => x"84808081",
   664 => x"842d8480",
   665 => x"8095d704",
   666 => x"9fe5c20b",
   667 => x"84808080",
   668 => x"b02d5473",
   669 => x"80d52e09",
   670 => x"810680db",
   671 => x"389fe5c3",
   672 => x"0b848080",
   673 => x"80b02d54",
   674 => x"7381aa2e",
   675 => x"09810680",
   676 => x"c638800b",
   677 => x"9fe1c40b",
   678 => x"84808080",
   679 => x"b02d5654",
   680 => x"7481e92e",
   681 => x"83388154",
   682 => x"7481eb2e",
   683 => x"8c388055",
   684 => x"73752e09",
   685 => x"810683b5",
   686 => x"389fe1cf",
   687 => x"0b848080",
   688 => x"80b02d55",
   689 => x"7491389f",
   690 => x"e1d00b84",
   691 => x"808080b0",
   692 => x"2d547382",
   693 => x"2e893880",
   694 => x"55848080",
   695 => x"98ed049f",
   696 => x"e1d10b84",
   697 => x"808080b0",
   698 => x"2d709fe5",
   699 => x"f40cff05",
   700 => x"9fe5e80c",
   701 => x"9fe1d20b",
   702 => x"84808080",
   703 => x"b02d9fe1",
   704 => x"d30b8480",
   705 => x"8080b02d",
   706 => x"58760577",
   707 => x"82802905",
   708 => x"709fe5dc",
   709 => x"0c9fe1d4",
   710 => x"0b848080",
   711 => x"80b02d70",
   712 => x"9fe5d40c",
   713 => x"9fe5ec08",
   714 => x"59575876",
   715 => x"802e81d7",
   716 => x"38885384",
   717 => x"8080a1ac",
   718 => x"529fe296",
   719 => x"51848080",
   720 => x"90c72d9f",
   721 => x"e0800882",
   722 => x"a4389fe5",
   723 => x"f4087084",
   724 => x"2b9fe5c4",
   725 => x"0c709fe5",
   726 => x"f00c9fe1",
   727 => x"e90b8480",
   728 => x"8080b02d",
   729 => x"9fe1e80b",
   730 => x"84808080",
   731 => x"b02d7182",
   732 => x"8029059f",
   733 => x"e1ea0b84",
   734 => x"808080b0",
   735 => x"2d708480",
   736 => x"8029129f",
   737 => x"e1eb0b84",
   738 => x"808080b0",
   739 => x"2d708180",
   740 => x"0a291270",
   741 => x"9fe1bc0c",
   742 => x"9fe5d408",
   743 => x"71299fe5",
   744 => x"dc080570",
   745 => x"9fe5fc0c",
   746 => x"9fe1f10b",
   747 => x"84808080",
   748 => x"b02d9fe1",
   749 => x"f00b8480",
   750 => x"8080b02d",
   751 => x"71828029",
   752 => x"059fe1f2",
   753 => x"0b848080",
   754 => x"80b02d70",
   755 => x"84808029",
   756 => x"129fe1f3",
   757 => x"0b848080",
   758 => x"80b02d70",
   759 => x"982b81f0",
   760 => x"0a067205",
   761 => x"709fe1c0",
   762 => x"0cfe117e",
   763 => x"2977059f",
   764 => x"e5e40c52",
   765 => x"59524354",
   766 => x"5e515259",
   767 => x"525d5759",
   768 => x"57848080",
   769 => x"98eb049f",
   770 => x"e1d60b84",
   771 => x"808080b0",
   772 => x"2d9fe1d5",
   773 => x"0b848080",
   774 => x"80b02d71",
   775 => x"82802905",
   776 => x"709fe5c4",
   777 => x"0c70a029",
   778 => x"83ff0570",
   779 => x"892a709f",
   780 => x"e5f00c9f",
   781 => x"e1db0b84",
   782 => x"808080b0",
   783 => x"2d9fe1da",
   784 => x"0b848080",
   785 => x"80b02d71",
   786 => x"82802905",
   787 => x"709fe1bc",
   788 => x"0c7b7129",
   789 => x"1e709fe5",
   790 => x"e40c7d9f",
   791 => x"e1c00c73",
   792 => x"059fe5fc",
   793 => x"0c555e51",
   794 => x"51555581",
   795 => x"55749fe0",
   796 => x"800c02a8",
   797 => x"050d0402",
   798 => x"ec050d76",
   799 => x"70872c71",
   800 => x"80ff0657",
   801 => x"55539fe5",
   802 => x"ec088a38",
   803 => x"72882c73",
   804 => x"81ff0656",
   805 => x"54739fe5",
   806 => x"d8082ea4",
   807 => x"389fe1c4",
   808 => x"529fe5dc",
   809 => x"08145184",
   810 => x"80808ea3",
   811 => x"2d9fe080",
   812 => x"08539fe0",
   813 => x"8008802e",
   814 => x"80c93873",
   815 => x"9fe5d80c",
   816 => x"9fe5ec08",
   817 => x"802ea038",
   818 => x"7484299f",
   819 => x"e1c40570",
   820 => x"08525384",
   821 => x"808083ec",
   822 => x"2d9fe080",
   823 => x"08f00a06",
   824 => x"55848080",
   825 => x"9a810474",
   826 => x"109fe1c4",
   827 => x"05708480",
   828 => x"80809b2d",
   829 => x"52538480",
   830 => x"80849d2d",
   831 => x"9fe08008",
   832 => x"55745372",
   833 => x"9fe0800c",
   834 => x"0294050d",
   835 => x"0402cc05",
   836 => x"0d7e605e",
   837 => x"5b8056ff",
   838 => x"0b9fe5d8",
   839 => x"0c9fe1c0",
   840 => x"089fe5e4",
   841 => x"0856579f",
   842 => x"e5ec0876",
   843 => x"2e8e389f",
   844 => x"e5f40884",
   845 => x"2b598480",
   846 => x"809ac304",
   847 => x"9fe5f008",
   848 => x"842b5980",
   849 => x"5a797927",
   850 => x"81e83879",
   851 => x"8f06a017",
   852 => x"575473a2",
   853 => x"38745284",
   854 => x"8080a2e4",
   855 => x"51848080",
   856 => x"81842d9f",
   857 => x"e1c45274",
   858 => x"51811555",
   859 => x"8480808e",
   860 => x"a32d9fe1",
   861 => x"c4568076",
   862 => x"84808080",
   863 => x"b02d5558",
   864 => x"73782e83",
   865 => x"38815873",
   866 => x"81e52e81",
   867 => x"9c388170",
   868 => x"7906555c",
   869 => x"73802e81",
   870 => x"90388b16",
   871 => x"84808080",
   872 => x"b02d9806",
   873 => x"58778181",
   874 => x"388b537c",
   875 => x"52755184",
   876 => x"808090c7",
   877 => x"2d9fe080",
   878 => x"0880ee38",
   879 => x"9c160851",
   880 => x"84808083",
   881 => x"ec2d9fe0",
   882 => x"8008841c",
   883 => x"0c9a1684",
   884 => x"8080809b",
   885 => x"2d518480",
   886 => x"80849d2d",
   887 => x"9fe08008",
   888 => x"9fe08008",
   889 => x"55559fe5",
   890 => x"ec08802e",
   891 => x"9f389416",
   892 => x"84808080",
   893 => x"9b2d5184",
   894 => x"8080849d",
   895 => x"2d9fe080",
   896 => x"08902b83",
   897 => x"fff00a06",
   898 => x"70165154",
   899 => x"73881c0c",
   900 => x"777b0c7c",
   901 => x"52848080",
   902 => x"a3845184",
   903 => x"80808184",
   904 => x"2d7b5484",
   905 => x"80809cff",
   906 => x"04811a5a",
   907 => x"8480809a",
   908 => x"c5049fe5",
   909 => x"ec08802e",
   910 => x"80c33876",
   911 => x"51848080",
   912 => x"98f72d9f",
   913 => x"e080089f",
   914 => x"e0800853",
   915 => x"848080a3",
   916 => x"98525784",
   917 => x"80808184",
   918 => x"2d7680ff",
   919 => x"fffff806",
   920 => x"547380ff",
   921 => x"fffff82e",
   922 => x"9438fe17",
   923 => x"9fe5f408",
   924 => x"299fe5fc",
   925 => x"08055584",
   926 => x"80809ac3",
   927 => x"04805473",
   928 => x"9fe0800c",
   929 => x"02b4050d",
   930 => x"0402e405",
   931 => x"0d787a71",
   932 => x"549fe5c8",
   933 => x"53555584",
   934 => x"80809a8d",
   935 => x"2d9fe080",
   936 => x"0881ff06",
   937 => x"5372802e",
   938 => x"80fe3884",
   939 => x"8080a3b0",
   940 => x"51848080",
   941 => x"85a92d9f",
   942 => x"e5cc0883",
   943 => x"ff05892a",
   944 => x"57807056",
   945 => x"56757725",
   946 => x"80fd389f",
   947 => x"e5d008fe",
   948 => x"059fe5f4",
   949 => x"08299fe5",
   950 => x"fc081176",
   951 => x"9fe5e808",
   952 => x"06057554",
   953 => x"52538480",
   954 => x"808ea32d",
   955 => x"9fe08008",
   956 => x"802e80c8",
   957 => x"38811570",
   958 => x"9fe5e808",
   959 => x"06545572",
   960 => x"94389fe5",
   961 => x"d0085184",
   962 => x"808098f7",
   963 => x"2d9fe080",
   964 => x"089fe5d0",
   965 => x"0c848014",
   966 => x"81175754",
   967 => x"767624ff",
   968 => x"aa388480",
   969 => x"809ec704",
   970 => x"74528480",
   971 => x"80a3cc51",
   972 => x"84808081",
   973 => x"842d8480",
   974 => x"809ec904",
   975 => x"9fe08008",
   976 => x"53848080",
   977 => x"9ec90481",
   978 => x"53729fe0",
   979 => x"800c029c",
   980 => x"050d049f",
   981 => x"e08c0802",
   982 => x"9fe08c0c",
   983 => x"ff3d0d80",
   984 => x"0b9fe08c",
   985 => x"08fc050c",
   986 => x"9fe08c08",
   987 => x"88050881",
   988 => x"06ff1170",
   989 => x"09709fe0",
   990 => x"8c088c05",
   991 => x"08069fe0",
   992 => x"8c08fc05",
   993 => x"08119fe0",
   994 => x"8c08fc05",
   995 => x"0c9fe08c",
   996 => x"08880508",
   997 => x"812a9fe0",
   998 => x"8c088805",
   999 => x"0c9fe08c",
  1000 => x"088c0508",
  1001 => x"109fe08c",
  1002 => x"088c050c",
  1003 => x"51515151",
  1004 => x"9fe08c08",
  1005 => x"88050880",
  1006 => x"2e8438ff",
  1007 => x"ab399fe0",
  1008 => x"8c08fc05",
  1009 => x"08709fe0",
  1010 => x"800c5183",
  1011 => x"3d0d9fe0",
  1012 => x"8c0c0400",
  1013 => x"00ffffff",
  1014 => x"ff00ffff",
  1015 => x"ffff00ff",
  1016 => x"ffffff00",
  1017 => x"436d645f",
  1018 => x"696e6974",
  1019 => x"0a000000",
  1020 => x"496e6974",
  1021 => x"69616c69",
  1022 => x"7a696e67",
  1023 => x"20534420",
  1024 => x"63617264",
  1025 => x"0a000000",
  1026 => x"48756e74",
  1027 => x"696e6720",
  1028 => x"666f7220",
  1029 => x"70617274",
  1030 => x"6974696f",
  1031 => x"6e0a0000",
  1032 => x"4f53445a",
  1033 => x"50553031",
  1034 => x"53595300",
  1035 => x"43616e27",
  1036 => x"74206c6f",
  1037 => x"61642066",
  1038 => x"69726d77",
  1039 => x"6172650a",
  1040 => x"00000000",
  1041 => x"4661696c",
  1042 => x"65642074",
  1043 => x"6f20696e",
  1044 => x"69746961",
  1045 => x"6c697a65",
  1046 => x"20534420",
  1047 => x"63617264",
  1048 => x"0a000000",
  1049 => x"52656164",
  1050 => x"696e6720",
  1051 => x"4d42520a",
  1052 => x"00000000",
  1053 => x"52656164",
  1054 => x"206f6620",
  1055 => x"4d425220",
  1056 => x"6661696c",
  1057 => x"65640a00",
  1058 => x"4d425220",
  1059 => x"73756363",
  1060 => x"65737366",
  1061 => x"756c6c79",
  1062 => x"20726561",
  1063 => x"640a0000",
  1064 => x"46415431",
  1065 => x"36202020",
  1066 => x"00000000",
  1067 => x"46415433",
  1068 => x"32202020",
  1069 => x"00000000",
  1070 => x"50617274",
  1071 => x"6974696f",
  1072 => x"6e636f75",
  1073 => x"6e742025",
  1074 => x"640a0000",
  1075 => x"4e6f2070",
  1076 => x"61727469",
  1077 => x"74696f6e",
  1078 => x"20736967",
  1079 => x"6e617475",
  1080 => x"72652066",
  1081 => x"6f756e64",
  1082 => x"0a000000",
  1083 => x"52656164",
  1084 => x"696e6720",
  1085 => x"626f6f74",
  1086 => x"20736563",
  1087 => x"746f7220",
  1088 => x"25640a00",
  1089 => x"52656164",
  1090 => x"20626f6f",
  1091 => x"74207365",
  1092 => x"63746f72",
  1093 => x"2066726f",
  1094 => x"6d206669",
  1095 => x"72737420",
  1096 => x"70617274",
  1097 => x"6974696f",
  1098 => x"6e0a0000",
  1099 => x"48756e74",
  1100 => x"696e6720",
  1101 => x"666f7220",
  1102 => x"66696c65",
  1103 => x"73797374",
  1104 => x"656d0a00",
  1105 => x"556e7375",
  1106 => x"70706f72",
  1107 => x"74656420",
  1108 => x"70617274",
  1109 => x"6974696f",
  1110 => x"6e207479",
  1111 => x"7065210d",
  1112 => x"00000000",
  1113 => x"52656164",
  1114 => x"696e6720",
  1115 => x"64697265",
  1116 => x"63746f72",
  1117 => x"79207365",
  1118 => x"63746f72",
  1119 => x"2025640a",
  1120 => x"00000000",
  1121 => x"66696c65",
  1122 => x"20222573",
  1123 => x"2220666f",
  1124 => x"756e640d",
  1125 => x"00000000",
  1126 => x"47657446",
  1127 => x"41544c69",
  1128 => x"6e6b2072",
  1129 => x"65747572",
  1130 => x"6e656420",
  1131 => x"25640a00",
  1132 => x"4f70656e",
  1133 => x"65642066",
  1134 => x"696c652c",
  1135 => x"206c6f61",
  1136 => x"64696e67",
  1137 => x"2e2e2e0a",
  1138 => x"00000000",
  1139 => x"43616e27",
  1140 => x"74206f70",
  1141 => x"656e2025",
  1142 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

