-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity DiagROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end DiagROM_ROM;

architecture arch of DiagROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ee040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"88080d80",
     5 => x"04848080",
     6 => x"80950471",
     7 => x"fd060872",
     8 => x"83060981",
     9 => x"05820583",
    10 => x"2b2a83ff",
    11 => x"ff065204",
    12 => x"71fc0608",
    13 => x"72830609",
    14 => x"81058305",
    15 => x"1010102a",
    16 => x"81ff0652",
    17 => x"0471fc06",
    18 => x"08848080",
    19 => x"a3cc7383",
    20 => x"06101005",
    21 => x"08067381",
    22 => x"ff067383",
    23 => x"06098105",
    24 => x"83051010",
    25 => x"102b0772",
    26 => x"fc060c51",
    27 => x"51040284",
    28 => x"05848080",
    29 => x"80880c84",
    30 => x"80808095",
    31 => x"0b848080",
    32 => x"93ce0400",
    33 => x"02c4050d",
    34 => x"0280c005",
    35 => x"9fe0e05b",
    36 => x"56807670",
    37 => x"84055808",
    38 => x"715e5e57",
    39 => x"7c708405",
    40 => x"5e085880",
    41 => x"5b77982a",
    42 => x"78882b59",
    43 => x"54738938",
    44 => x"765e8480",
    45 => x"8083e204",
    46 => x"7b802e81",
    47 => x"fd38805c",
    48 => x"7380e42e",
    49 => x"a1387380",
    50 => x"e4268e38",
    51 => x"7380e32e",
    52 => x"819a3884",
    53 => x"808082fa",
    54 => x"047380f3",
    55 => x"2e80f538",
    56 => x"84808082",
    57 => x"fa047584",
    58 => x"1771087e",
    59 => x"5c555752",
    60 => x"7280258e",
    61 => x"38ad5184",
    62 => x"808092fb",
    63 => x"2d720981",
    64 => x"05537280",
    65 => x"2ebe3887",
    66 => x"55729c2a",
    67 => x"73842b54",
    68 => x"5271802e",
    69 => x"83388159",
    70 => x"8972258a",
    71 => x"38b71252",
    72 => x"84808082",
    73 => x"a904b012",
    74 => x"5278802e",
    75 => x"89387151",
    76 => x"84808092",
    77 => x"fb2dff15",
    78 => x"55748025",
    79 => x"cc388480",
    80 => x"8082cc04",
    81 => x"b0518480",
    82 => x"8092fb2d",
    83 => x"80538480",
    84 => x"80839304",
    85 => x"75841771",
    86 => x"0870545c",
    87 => x"57528480",
    88 => x"80938f2d",
    89 => x"7b538480",
    90 => x"80839304",
    91 => x"75841771",
    92 => x"08565752",
    93 => x"84808083",
    94 => x"ca04a551",
    95 => x"84808092",
    96 => x"fb2d7351",
    97 => x"84808092",
    98 => x"fb2d8217",
    99 => x"57848080",
   100 => x"83d50472",
   101 => x"ff145452",
   102 => x"807225b9",
   103 => x"38797081",
   104 => x"055b8480",
   105 => x"8080b02d",
   106 => x"70525484",
   107 => x"808092fb",
   108 => x"2d811757",
   109 => x"84808083",
   110 => x"930473a5",
   111 => x"2e098106",
   112 => x"8938815c",
   113 => x"84808083",
   114 => x"d5047351",
   115 => x"84808092",
   116 => x"fb2d8117",
   117 => x"57811b5b",
   118 => x"837b25fd",
   119 => x"c83873fd",
   120 => x"bb387d9f",
   121 => x"e0800c02",
   122 => x"bc050d04",
   123 => x"02f4050d",
   124 => x"7470882a",
   125 => x"83fe8006",
   126 => x"7072982a",
   127 => x"0772882b",
   128 => x"87fc8080",
   129 => x"0673982b",
   130 => x"81f00a06",
   131 => x"71730707",
   132 => x"9fe0800c",
   133 => x"56515351",
   134 => x"028c050d",
   135 => x"0402f805",
   136 => x"0d73882b",
   137 => x"83fe8006",
   138 => x"0284058e",
   139 => x"05848080",
   140 => x"80b02d71",
   141 => x"079fe080",
   142 => x"0c510288",
   143 => x"050d0402",
   144 => x"f8050d73",
   145 => x"70902b71",
   146 => x"902a079f",
   147 => x"e0800c52",
   148 => x"0288050d",
   149 => x"0402f805",
   150 => x"0d735170",
   151 => x"802e8c38",
   152 => x"709fe1a0",
   153 => x"0c800b9f",
   154 => x"e1a80c9f",
   155 => x"e1a80852",
   156 => x"7198389f",
   157 => x"e1a00884",
   158 => x"119fe1a0",
   159 => x"0c70089f",
   160 => x"e1a40c51",
   161 => x"84808085",
   162 => x"94049fe1",
   163 => x"a408882b",
   164 => x"9fe1a40c",
   165 => x"81128306",
   166 => x"9fe1a80c",
   167 => x"9fe1a408",
   168 => x"982c9fe0",
   169 => x"800c0288",
   170 => x"050d0402",
   171 => x"e8050d77",
   172 => x"70525684",
   173 => x"808084d5",
   174 => x"2d9fe080",
   175 => x"08528053",
   176 => x"71802e97",
   177 => x"38811353",
   178 => x"80518480",
   179 => x"8084d52d",
   180 => x"9fe08008",
   181 => x"52848080",
   182 => x"85c00482",
   183 => x"13548155",
   184 => x"900b86e9",
   185 => x"808423a0",
   186 => x"810b86e9",
   187 => x"80802386",
   188 => x"e9808022",
   189 => x"52800b86",
   190 => x"e9808023",
   191 => x"86e98080",
   192 => x"2253800b",
   193 => x"86e98080",
   194 => x"2386e980",
   195 => x"80227083",
   196 => x"ffff0673",
   197 => x"882a7081",
   198 => x"06515451",
   199 => x"5371802e",
   200 => x"81a43874",
   201 => x"802e80e0",
   202 => x"38728280",
   203 => x"862e0981",
   204 => x"06819338",
   205 => x"8055fed5",
   206 => x"ca0b86e9",
   207 => x"80802386",
   208 => x"e9808022",
   209 => x"52810b86",
   210 => x"e9808023",
   211 => x"86e98080",
   212 => x"22527486",
   213 => x"e9808023",
   214 => x"86e98080",
   215 => x"22527386",
   216 => x"e9808023",
   217 => x"86e98080",
   218 => x"22527486",
   219 => x"e9808023",
   220 => x"86e98080",
   221 => x"22527486",
   222 => x"e9808023",
   223 => x"86e98080",
   224 => x"22528480",
   225 => x"8087c604",
   226 => x"73812a82",
   227 => x"80800752",
   228 => x"72722e09",
   229 => x"8106af38",
   230 => x"75518480",
   231 => x"8084d52d",
   232 => x"9fe08008",
   233 => x"53ff1454",
   234 => x"73ff2ea7",
   235 => x"387286e9",
   236 => x"80803486",
   237 => x"e9808033",
   238 => x"5272802e",
   239 => x"e8388051",
   240 => x"84808087",
   241 => x"9a04910b",
   242 => x"86e98084",
   243 => x"23848080",
   244 => x"85e00491",
   245 => x"0b86e980",
   246 => x"8423810b",
   247 => x"9fe0800c",
   248 => x"0298050d",
   249 => x"0402f405",
   250 => x"0d86e980",
   251 => x"8152ff72",
   252 => x"34713353",
   253 => x"ff723472",
   254 => x"882b83fe",
   255 => x"80067233",
   256 => x"7081ff06",
   257 => x"515253ff",
   258 => x"72347271",
   259 => x"07882b72",
   260 => x"337081ff",
   261 => x"06515253",
   262 => x"ff723472",
   263 => x"7107882b",
   264 => x"72337081",
   265 => x"ff067207",
   266 => x"9fe0800c",
   267 => x"5253028c",
   268 => x"050d0402",
   269 => x"ec050d76",
   270 => x"78848080",
   271 => x"a3dc5355",
   272 => x"55848080",
   273 => x"938f2d74",
   274 => x"86e98081",
   275 => x"34848080",
   276 => x"a3ec5184",
   277 => x"8080938f",
   278 => x"2d9fe1ac",
   279 => x"08853873",
   280 => x"892b5484",
   281 => x"8080a3fc",
   282 => x"51848080",
   283 => x"938f2d73",
   284 => x"982a5372",
   285 => x"86e98081",
   286 => x"34848080",
   287 => x"a48c5184",
   288 => x"8080938f",
   289 => x"2d73902a",
   290 => x"537286e9",
   291 => x"80813484",
   292 => x"8080a49c",
   293 => x"51848080",
   294 => x"938f2d73",
   295 => x"882a5372",
   296 => x"86e98081",
   297 => x"34848080",
   298 => x"a4ac5184",
   299 => x"8080938f",
   300 => x"2d7386e9",
   301 => x"80813484",
   302 => x"8080a4bc",
   303 => x"51848080",
   304 => x"938f2d84",
   305 => x"8080a4cc",
   306 => x"51848080",
   307 => x"938f2d74",
   308 => x"902a5372",
   309 => x"86e98081",
   310 => x"3486e980",
   311 => x"81337081",
   312 => x"ff065153",
   313 => x"82b8bf54",
   314 => x"7281ff2e",
   315 => x"09810699",
   316 => x"38ff0b86",
   317 => x"e9808134",
   318 => x"86e98081",
   319 => x"337081ff",
   320 => x"06ff1656",
   321 => x"515373e0",
   322 => x"3872842a",
   323 => x"b0055184",
   324 => x"808092fb",
   325 => x"2d72bf06",
   326 => x"b0075184",
   327 => x"808092fb",
   328 => x"2d725284",
   329 => x"8080a4e4",
   330 => x"51848080",
   331 => x"81842d72",
   332 => x"9fe0800c",
   333 => x"0294050d",
   334 => x"0402fc05",
   335 => x"0d81c751",
   336 => x"ff0b86e9",
   337 => x"808134ff",
   338 => x"11517080",
   339 => x"25f23802",
   340 => x"84050d04",
   341 => x"02f0050d",
   342 => x"8480808a",
   343 => x"b92d819c",
   344 => x"9f538052",
   345 => x"87fc80f7",
   346 => x"51848080",
   347 => x"88b32d9f",
   348 => x"e0800854",
   349 => x"9fe08008",
   350 => x"812e0981",
   351 => x"0680ea38",
   352 => x"9fe08008",
   353 => x"52848080",
   354 => x"a4f45184",
   355 => x"80808184",
   356 => x"2dff0b86",
   357 => x"e9808134",
   358 => x"820a5284",
   359 => x"9c80e951",
   360 => x"84808088",
   361 => x"b32d9fe0",
   362 => x"8008a138",
   363 => x"9fe08008",
   364 => x"52848080",
   365 => x"a5805184",
   366 => x"80808184",
   367 => x"2dff0b86",
   368 => x"e9808134",
   369 => x"73538480",
   370 => x"808c8104",
   371 => x"9fe08008",
   372 => x"52848080",
   373 => x"a5805184",
   374 => x"80808184",
   375 => x"2d848080",
   376 => x"8ab92d84",
   377 => x"80808bfa",
   378 => x"049fe080",
   379 => x"08528480",
   380 => x"80a4f451",
   381 => x"84808081",
   382 => x"842dff13",
   383 => x"5372fee2",
   384 => x"38729fe0",
   385 => x"800c0290",
   386 => x"050d0402",
   387 => x"f4050dff",
   388 => x"0b86e980",
   389 => x"81348480",
   390 => x"80a58c51",
   391 => x"84808093",
   392 => x"8f2d9353",
   393 => x"805287fc",
   394 => x"80c15184",
   395 => x"808088b3",
   396 => x"2d9fe080",
   397 => x"08a1389f",
   398 => x"e0800852",
   399 => x"848080a5",
   400 => x"98518480",
   401 => x"8081842d",
   402 => x"ff0b86e9",
   403 => x"80813481",
   404 => x"53848080",
   405 => x"8cf5049f",
   406 => x"e0800852",
   407 => x"848080a5",
   408 => x"98518480",
   409 => x"8081842d",
   410 => x"8480808a",
   411 => x"b92dff13",
   412 => x"5372ffb0",
   413 => x"38729fe0",
   414 => x"800c028c",
   415 => x"050d0402",
   416 => x"f0050d84",
   417 => x"80808ab9",
   418 => x"2d83aa52",
   419 => x"849c80c8",
   420 => x"51848080",
   421 => x"88b32d9f",
   422 => x"e080089f",
   423 => x"e0800853",
   424 => x"848080a5",
   425 => x"a4525384",
   426 => x"80808184",
   427 => x"2d72812e",
   428 => x"098106a7",
   429 => x"38848080",
   430 => x"87e52d9f",
   431 => x"e0800883",
   432 => x"ffff0653",
   433 => x"7283aa2e",
   434 => x"ba389fe0",
   435 => x"80085284",
   436 => x"8080a5bc",
   437 => x"51848080",
   438 => x"81842d84",
   439 => x"80808c8b",
   440 => x"2d848080",
   441 => x"8dfb0481",
   442 => x"54848080",
   443 => x"8fb10484",
   444 => x"8080a5d4",
   445 => x"51848080",
   446 => x"81842d80",
   447 => x"54848080",
   448 => x"8fb104ff",
   449 => x"0b86e980",
   450 => x"8134b153",
   451 => x"8480808a",
   452 => x"d42d9fe0",
   453 => x"8008802e",
   454 => x"81883880",
   455 => x"5287fc80",
   456 => x"fa518480",
   457 => x"8088b32d",
   458 => x"9fe08008",
   459 => x"80e3389f",
   460 => x"e0800852",
   461 => x"848080a5",
   462 => x"f0518480",
   463 => x"8081842d",
   464 => x"ff0b86e9",
   465 => x"80813486",
   466 => x"e9808133",
   467 => x"7081ff06",
   468 => x"70548480",
   469 => x"80a5fc53",
   470 => x"51538480",
   471 => x"8081842d",
   472 => x"ff0b86e9",
   473 => x"808134ff",
   474 => x"0b86e980",
   475 => x"8134ff0b",
   476 => x"86e98081",
   477 => x"34ff0b86",
   478 => x"e9808134",
   479 => x"72862a70",
   480 => x"81067056",
   481 => x"51537280",
   482 => x"2ea73884",
   483 => x"80808de7",
   484 => x"049fe080",
   485 => x"08528480",
   486 => x"80a5f051",
   487 => x"84808081",
   488 => x"842d7282",
   489 => x"2efec838",
   490 => x"ff135372",
   491 => x"fede3872",
   492 => x"54739fe0",
   493 => x"800c0290",
   494 => x"050d0402",
   495 => x"f4050d81",
   496 => x"0b9fe1ac",
   497 => x"0ca00b86",
   498 => x"e9808934",
   499 => x"830b86e9",
   500 => x"80853484",
   501 => x"80808ab9",
   502 => x"2d848080",
   503 => x"a68c5184",
   504 => x"8080938f",
   505 => x"2d820b86",
   506 => x"e9808534",
   507 => x"87538052",
   508 => x"84d480c0",
   509 => x"51848080",
   510 => x"88b32d9f",
   511 => x"e0800881",
   512 => x"2e098106",
   513 => x"86389fe0",
   514 => x"80085384",
   515 => x"8080a69c",
   516 => x"51848080",
   517 => x"938f2d72",
   518 => x"822e0981",
   519 => x"06953884",
   520 => x"8080a6b0",
   521 => x"51848080",
   522 => x"938f2d80",
   523 => x"53848080",
   524 => x"91a404ff",
   525 => x"135372ff",
   526 => x"b5388480",
   527 => x"80a6d051",
   528 => x"84808093",
   529 => x"8f2d8480",
   530 => x"808cff2d",
   531 => x"9fe08008",
   532 => x"9fe1ac0c",
   533 => x"9fe08008",
   534 => x"802e8d38",
   535 => x"848080a6",
   536 => x"ec518480",
   537 => x"80938f2d",
   538 => x"848080a7",
   539 => x"80518480",
   540 => x"80938f2d",
   541 => x"815287fc",
   542 => x"80d05184",
   543 => x"808088b3",
   544 => x"2dff0b86",
   545 => x"e9808134",
   546 => x"830b86e9",
   547 => x"808534ff",
   548 => x"0b86e980",
   549 => x"81348480",
   550 => x"80a79051",
   551 => x"84808093",
   552 => x"8f2d8153",
   553 => x"729fe080",
   554 => x"0c028c05",
   555 => x"0d04800b",
   556 => x"9fe0800c",
   557 => x"0402e405",
   558 => x"0d787a57",
   559 => x"54807654",
   560 => x"74538480",
   561 => x"80a79c52",
   562 => x"57848080",
   563 => x"81842dff",
   564 => x"0b86e980",
   565 => x"8134820b",
   566 => x"86e98085",
   567 => x"34810b86",
   568 => x"e9808934",
   569 => x"ff0b86e9",
   570 => x"80813473",
   571 => x"5287fc80",
   572 => x"d1518480",
   573 => x"8088b32d",
   574 => x"80dbc6df",
   575 => x"559fe080",
   576 => x"08772e9a",
   577 => x"389fe080",
   578 => x"08537352",
   579 => x"848080a7",
   580 => x"b4518480",
   581 => x"8081842d",
   582 => x"84808092",
   583 => x"f104ff0b",
   584 => x"86e98081",
   585 => x"3486e980",
   586 => x"81337081",
   587 => x"ff065154",
   588 => x"7381fe2e",
   589 => x"098106a4",
   590 => x"3880ff54",
   591 => x"84808087",
   592 => x"e52d9fe0",
   593 => x"80087670",
   594 => x"8405580c",
   595 => x"ff145473",
   596 => x"8025e938",
   597 => x"81578480",
   598 => x"8092e304",
   599 => x"ff155574",
   600 => x"ffbc38ff",
   601 => x"0b86e980",
   602 => x"8134830b",
   603 => x"86e98085",
   604 => x"34769fe0",
   605 => x"800c029c",
   606 => x"050d0402",
   607 => x"fc050d72",
   608 => x"7086ea80",
   609 => x"800c9fe0",
   610 => x"800c0284",
   611 => x"050d0402",
   612 => x"ec050d80",
   613 => x"77565474",
   614 => x"70840556",
   615 => x"08518053",
   616 => x"70982a71",
   617 => x"882b5252",
   618 => x"71802e98",
   619 => x"387186ea",
   620 => x"80800c81",
   621 => x"14811454",
   622 => x"54837325",
   623 => x"e3388480",
   624 => x"80939704",
   625 => x"739fe080",
   626 => x"0c029405",
   627 => x"0d0402f8",
   628 => x"050d8480",
   629 => x"80a7d451",
   630 => x"84808093",
   631 => x"8f2d8480",
   632 => x"808fbb2d",
   633 => x"9fe08008",
   634 => x"802ebb38",
   635 => x"848080a7",
   636 => x"ec518480",
   637 => x"80938f2d",
   638 => x"84808095",
   639 => x"882d8052",
   640 => x"848080a8",
   641 => x"84518480",
   642 => x"80a0ff2d",
   643 => x"9fe08008",
   644 => x"802e8738",
   645 => x"84808080",
   646 => x"8c2d8480",
   647 => x"80a89051",
   648 => x"84808093",
   649 => x"8f2d8480",
   650 => x"80a8a851",
   651 => x"84808093",
   652 => x"8f2d800b",
   653 => x"9fe0800c",
   654 => x"0288050d",
   655 => x"0402e805",
   656 => x"0d77797b",
   657 => x"58555580",
   658 => x"53727625",
   659 => x"af387470",
   660 => x"81055684",
   661 => x"808080b0",
   662 => x"2d747081",
   663 => x"05568480",
   664 => x"8080b02d",
   665 => x"52527171",
   666 => x"2e893881",
   667 => x"51848080",
   668 => x"94fe0481",
   669 => x"13538480",
   670 => x"8094c904",
   671 => x"8051709f",
   672 => x"e0800c02",
   673 => x"98050d04",
   674 => x"02d8050d",
   675 => x"ff0b9fe5",
   676 => x"d80c800b",
   677 => x"9fe5ec0c",
   678 => x"848080a8",
   679 => x"c8518480",
   680 => x"80938f2d",
   681 => x"9fe1c452",
   682 => x"80518480",
   683 => x"8091b52d",
   684 => x"9fe08008",
   685 => x"549fe080",
   686 => x"08953884",
   687 => x"8080a8d8",
   688 => x"51848080",
   689 => x"938f2d73",
   690 => x"55848080",
   691 => x"9ce30484",
   692 => x"8080a8ec",
   693 => x"51848080",
   694 => x"938f2d80",
   695 => x"56810b9f",
   696 => x"e1b80c88",
   697 => x"53848080",
   698 => x"a984529f",
   699 => x"e1fa5184",
   700 => x"808094bd",
   701 => x"2d9fe080",
   702 => x"08762e09",
   703 => x"81068938",
   704 => x"9fe08008",
   705 => x"9fe1b80c",
   706 => x"88538480",
   707 => x"80a99052",
   708 => x"9fe29651",
   709 => x"84808094",
   710 => x"bd2d9fe0",
   711 => x"80088938",
   712 => x"9fe08008",
   713 => x"9fe1b80c",
   714 => x"9fe1b808",
   715 => x"52848080",
   716 => x"a99c5184",
   717 => x"80808184",
   718 => x"2d9fe1b8",
   719 => x"08802e81",
   720 => x"c1389fe5",
   721 => x"8a0b8480",
   722 => x"8080b02d",
   723 => x"9fe58b0b",
   724 => x"84808080",
   725 => x"b02d7198",
   726 => x"2b71902b",
   727 => x"079fe58c",
   728 => x"0b848080",
   729 => x"80b02d70",
   730 => x"882b7207",
   731 => x"9fe58d0b",
   732 => x"84808080",
   733 => x"b02d7107",
   734 => x"9fe5c20b",
   735 => x"84808080",
   736 => x"b02d9fe5",
   737 => x"c30b8480",
   738 => x"8080b02d",
   739 => x"71882b07",
   740 => x"535f5452",
   741 => x"5a565755",
   742 => x"7381abaa",
   743 => x"2e098106",
   744 => x"94387551",
   745 => x"84808083",
   746 => x"ec2d9fe0",
   747 => x"80085684",
   748 => x"808097ce",
   749 => x"047382d4",
   750 => x"d52e9338",
   751 => x"848080a9",
   752 => x"b0518480",
   753 => x"80938f2d",
   754 => x"84808099",
   755 => x"cd047552",
   756 => x"848080a9",
   757 => x"d0518480",
   758 => x"8081842d",
   759 => x"9fe1c452",
   760 => x"75518480",
   761 => x"8091b52d",
   762 => x"9fe08008",
   763 => x"559fe080",
   764 => x"08802e84",
   765 => x"ee388480",
   766 => x"80a9e851",
   767 => x"84808093",
   768 => x"8f2d8480",
   769 => x"80aa9051",
   770 => x"84808081",
   771 => x"842d8853",
   772 => x"848080a9",
   773 => x"90529fe2",
   774 => x"96518480",
   775 => x"8094bd2d",
   776 => x"9fe08008",
   777 => x"8d38810b",
   778 => x"9fe5ec0c",
   779 => x"84808098",
   780 => x"de048853",
   781 => x"848080a9",
   782 => x"84529fe1",
   783 => x"fa518480",
   784 => x"8094bd2d",
   785 => x"9fe08008",
   786 => x"802e9338",
   787 => x"848080aa",
   788 => x"a8518480",
   789 => x"8081842d",
   790 => x"84808099",
   791 => x"cd049fe5",
   792 => x"c20b8480",
   793 => x"8080b02d",
   794 => x"547380d5",
   795 => x"2e098106",
   796 => x"80db389f",
   797 => x"e5c30b84",
   798 => x"808080b0",
   799 => x"2d547381",
   800 => x"aa2e0981",
   801 => x"0680c638",
   802 => x"800b9fe1",
   803 => x"c40b8480",
   804 => x"8080b02d",
   805 => x"56547481",
   806 => x"e92e8338",
   807 => x"81547481",
   808 => x"eb2e8c38",
   809 => x"80557375",
   810 => x"2e098106",
   811 => x"83b5389f",
   812 => x"e1cf0b84",
   813 => x"808080b0",
   814 => x"2d557491",
   815 => x"389fe1d0",
   816 => x"0b848080",
   817 => x"80b02d54",
   818 => x"73822e89",
   819 => x"38805584",
   820 => x"80809ce3",
   821 => x"049fe1d1",
   822 => x"0b848080",
   823 => x"80b02d70",
   824 => x"9fe5f40c",
   825 => x"ff059fe5",
   826 => x"e80c9fe1",
   827 => x"d20b8480",
   828 => x"8080b02d",
   829 => x"9fe1d30b",
   830 => x"84808080",
   831 => x"b02d5876",
   832 => x"05778280",
   833 => x"2905709f",
   834 => x"e5dc0c9f",
   835 => x"e1d40b84",
   836 => x"808080b0",
   837 => x"2d709fe5",
   838 => x"d40c9fe5",
   839 => x"ec085957",
   840 => x"5876802e",
   841 => x"81d73888",
   842 => x"53848080",
   843 => x"a990529f",
   844 => x"e2965184",
   845 => x"808094bd",
   846 => x"2d9fe080",
   847 => x"0882a438",
   848 => x"9fe5f408",
   849 => x"70842b9f",
   850 => x"e5c40c70",
   851 => x"9fe5f00c",
   852 => x"9fe1e90b",
   853 => x"84808080",
   854 => x"b02d9fe1",
   855 => x"e80b8480",
   856 => x"8080b02d",
   857 => x"71828029",
   858 => x"059fe1ea",
   859 => x"0b848080",
   860 => x"80b02d70",
   861 => x"84808029",
   862 => x"129fe1eb",
   863 => x"0b848080",
   864 => x"80b02d70",
   865 => x"81800a29",
   866 => x"12709fe1",
   867 => x"bc0c9fe5",
   868 => x"d4087129",
   869 => x"9fe5dc08",
   870 => x"05709fe5",
   871 => x"fc0c9fe1",
   872 => x"f10b8480",
   873 => x"8080b02d",
   874 => x"9fe1f00b",
   875 => x"84808080",
   876 => x"b02d7182",
   877 => x"8029059f",
   878 => x"e1f20b84",
   879 => x"808080b0",
   880 => x"2d708480",
   881 => x"8029129f",
   882 => x"e1f30b84",
   883 => x"808080b0",
   884 => x"2d70982b",
   885 => x"81f00a06",
   886 => x"7205709f",
   887 => x"e1c00cfe",
   888 => x"117e2977",
   889 => x"059fe5e4",
   890 => x"0c525952",
   891 => x"43545e51",
   892 => x"5259525d",
   893 => x"57595784",
   894 => x"80809ce1",
   895 => x"049fe1d6",
   896 => x"0b848080",
   897 => x"80b02d9f",
   898 => x"e1d50b84",
   899 => x"808080b0",
   900 => x"2d718280",
   901 => x"2905709f",
   902 => x"e5c40c70",
   903 => x"a02983ff",
   904 => x"0570892a",
   905 => x"709fe5f0",
   906 => x"0c9fe1db",
   907 => x"0b848080",
   908 => x"80b02d9f",
   909 => x"e1da0b84",
   910 => x"808080b0",
   911 => x"2d718280",
   912 => x"2905709f",
   913 => x"e1bc0c7b",
   914 => x"71291e70",
   915 => x"9fe5e40c",
   916 => x"7d9fe1c0",
   917 => x"0c73059f",
   918 => x"e5fc0c55",
   919 => x"5e515155",
   920 => x"55815574",
   921 => x"9fe0800c",
   922 => x"02a8050d",
   923 => x"0402ec05",
   924 => x"0d767087",
   925 => x"2c7180ff",
   926 => x"06575553",
   927 => x"9fe5ec08",
   928 => x"8a387288",
   929 => x"2c7381ff",
   930 => x"06565473",
   931 => x"9fe5d808",
   932 => x"2ea4389f",
   933 => x"e1c4529f",
   934 => x"e5dc0814",
   935 => x"51848080",
   936 => x"91b52d9f",
   937 => x"e0800853",
   938 => x"9fe08008",
   939 => x"802e80c9",
   940 => x"38739fe5",
   941 => x"d80c9fe5",
   942 => x"ec08802e",
   943 => x"a0387484",
   944 => x"299fe1c4",
   945 => x"05700852",
   946 => x"53848080",
   947 => x"83ec2d9f",
   948 => x"e08008f0",
   949 => x"0a065584",
   950 => x"80809df7",
   951 => x"0474109f",
   952 => x"e1c40570",
   953 => x"84808080",
   954 => x"9b2d5253",
   955 => x"84808084",
   956 => x"9d2d9fe0",
   957 => x"80085574",
   958 => x"53729fe0",
   959 => x"800c0294",
   960 => x"050d0402",
   961 => x"cc050d7e",
   962 => x"605e5b80",
   963 => x"56ff0b9f",
   964 => x"e5d80c9f",
   965 => x"e1c0089f",
   966 => x"e5e40856",
   967 => x"579fe5ec",
   968 => x"08762e8e",
   969 => x"389fe5f4",
   970 => x"08842b59",
   971 => x"8480809e",
   972 => x"b9049fe5",
   973 => x"f008842b",
   974 => x"59805a79",
   975 => x"792781e8",
   976 => x"38798f06",
   977 => x"a0175754",
   978 => x"73a23874",
   979 => x"52848080",
   980 => x"aac85184",
   981 => x"80808184",
   982 => x"2d9fe1c4",
   983 => x"52745181",
   984 => x"15558480",
   985 => x"8091b52d",
   986 => x"9fe1c456",
   987 => x"80768480",
   988 => x"8080b02d",
   989 => x"55587378",
   990 => x"2e833881",
   991 => x"587381e5",
   992 => x"2e819c38",
   993 => x"81707906",
   994 => x"555c7380",
   995 => x"2e819038",
   996 => x"8b168480",
   997 => x"8080b02d",
   998 => x"98065877",
   999 => x"8181388b",
  1000 => x"537c5275",
  1001 => x"51848080",
  1002 => x"94bd2d9f",
  1003 => x"e0800880",
  1004 => x"ee389c16",
  1005 => x"08518480",
  1006 => x"8083ec2d",
  1007 => x"9fe08008",
  1008 => x"841c0c9a",
  1009 => x"16848080",
  1010 => x"809b2d51",
  1011 => x"84808084",
  1012 => x"9d2d9fe0",
  1013 => x"80089fe0",
  1014 => x"80085555",
  1015 => x"9fe5ec08",
  1016 => x"802e9f38",
  1017 => x"94168480",
  1018 => x"80809b2d",
  1019 => x"51848080",
  1020 => x"849d2d9f",
  1021 => x"e0800890",
  1022 => x"2b83fff0",
  1023 => x"0a067016",
  1024 => x"51547388",
  1025 => x"1c0c777b",
  1026 => x"0c7c5284",
  1027 => x"8080aae8",
  1028 => x"51848080",
  1029 => x"81842d7b",
  1030 => x"54848080",
  1031 => x"a0f50481",
  1032 => x"1a5a8480",
  1033 => x"809ebb04",
  1034 => x"9fe5ec08",
  1035 => x"802e80c3",
  1036 => x"38765184",
  1037 => x"80809ced",
  1038 => x"2d9fe080",
  1039 => x"089fe080",
  1040 => x"08538480",
  1041 => x"80aafc52",
  1042 => x"57848080",
  1043 => x"81842d76",
  1044 => x"80ffffff",
  1045 => x"f8065473",
  1046 => x"80ffffff",
  1047 => x"f82e9438",
  1048 => x"fe179fe5",
  1049 => x"f408299f",
  1050 => x"e5fc0805",
  1051 => x"55848080",
  1052 => x"9eb90480",
  1053 => x"54739fe0",
  1054 => x"800c02b4",
  1055 => x"050d0402",
  1056 => x"e4050d78",
  1057 => x"7a71549f",
  1058 => x"e5c85355",
  1059 => x"55848080",
  1060 => x"9e832d9f",
  1061 => x"e0800881",
  1062 => x"ff065372",
  1063 => x"802e80fe",
  1064 => x"38848080",
  1065 => x"ab945184",
  1066 => x"8080938f",
  1067 => x"2d9fe5cc",
  1068 => x"0883ff05",
  1069 => x"892a5780",
  1070 => x"70565675",
  1071 => x"772580fd",
  1072 => x"389fe5d0",
  1073 => x"08fe059f",
  1074 => x"e5f40829",
  1075 => x"9fe5fc08",
  1076 => x"11769fe5",
  1077 => x"e8080605",
  1078 => x"75545253",
  1079 => x"84808091",
  1080 => x"b52d9fe0",
  1081 => x"8008802e",
  1082 => x"80c83881",
  1083 => x"15709fe5",
  1084 => x"e8080654",
  1085 => x"55729438",
  1086 => x"9fe5d008",
  1087 => x"51848080",
  1088 => x"9ced2d9f",
  1089 => x"e080089f",
  1090 => x"e5d00c84",
  1091 => x"80148117",
  1092 => x"57547676",
  1093 => x"24ffaa38",
  1094 => x"848080a2",
  1095 => x"bd047452",
  1096 => x"848080ab",
  1097 => x"b0518480",
  1098 => x"8081842d",
  1099 => x"848080a2",
  1100 => x"bf049fe0",
  1101 => x"80085384",
  1102 => x"8080a2bf",
  1103 => x"04815372",
  1104 => x"9fe0800c",
  1105 => x"029c050d",
  1106 => x"049fe08c",
  1107 => x"08029fe0",
  1108 => x"8c0cff3d",
  1109 => x"0d800b9f",
  1110 => x"e08c08fc",
  1111 => x"050c9fe0",
  1112 => x"8c088805",
  1113 => x"088106ff",
  1114 => x"11700970",
  1115 => x"9fe08c08",
  1116 => x"8c050806",
  1117 => x"9fe08c08",
  1118 => x"fc050811",
  1119 => x"9fe08c08",
  1120 => x"fc050c9f",
  1121 => x"e08c0888",
  1122 => x"0508812a",
  1123 => x"9fe08c08",
  1124 => x"88050c9f",
  1125 => x"e08c088c",
  1126 => x"0508109f",
  1127 => x"e08c088c",
  1128 => x"050c5151",
  1129 => x"51519fe0",
  1130 => x"8c088805",
  1131 => x"08802e84",
  1132 => x"38ffab39",
  1133 => x"9fe08c08",
  1134 => x"fc050870",
  1135 => x"9fe0800c",
  1136 => x"51833d0d",
  1137 => x"9fe08c0c",
  1138 => x"04000000",
  1139 => x"00ffffff",
  1140 => x"ff00ffff",
  1141 => x"ffff00ff",
  1142 => x"ffffff00",
  1143 => x"496e2063",
  1144 => x"6d645f77",
  1145 => x"72697465",
  1146 => x"0a000000",
  1147 => x"436f6d6d",
  1148 => x"616e6420",
  1149 => x"73656e74",
  1150 => x"0a000000",
  1151 => x"53656e64",
  1152 => x"696e6720",
  1153 => x"4c424121",
  1154 => x"0a000000",
  1155 => x"53656e74",
  1156 => x"20317374",
  1157 => x"20627974",
  1158 => x"650a0000",
  1159 => x"53656e74",
  1160 => x"20326e64",
  1161 => x"20627974",
  1162 => x"650a0000",
  1163 => x"53656e74",
  1164 => x"20337264",
  1165 => x"20627974",
  1166 => x"650a0000",
  1167 => x"53656e74",
  1168 => x"20347468",
  1169 => x"20627974",
  1170 => x"650a0000",
  1171 => x"53656e64",
  1172 => x"696e6720",
  1173 => x"43524320",
  1174 => x"2d206966",
  1175 => x"20616e79",
  1176 => x"0a000000",
  1177 => x"476f7420",
  1178 => x"72657375",
  1179 => x"6c742025",
  1180 => x"64200a00",
  1181 => x"434d4435",
  1182 => x"35202564",
  1183 => x"0a000000",
  1184 => x"434d4434",
  1185 => x"31202564",
  1186 => x"0a000000",
  1187 => x"436d645f",
  1188 => x"696e6974",
  1189 => x"0a000000",
  1190 => x"696e6974",
  1191 => x"2025640a",
  1192 => x"20200000",
  1193 => x"636d645f",
  1194 => x"434d4438",
  1195 => x"20726573",
  1196 => x"706f6e73",
  1197 => x"653a2025",
  1198 => x"640a0000",
  1199 => x"434d4438",
  1200 => x"5f342072",
  1201 => x"6573706f",
  1202 => x"6e73653a",
  1203 => x"2025640a",
  1204 => x"00000000",
  1205 => x"53444843",
  1206 => x"20496e69",
  1207 => x"7469616c",
  1208 => x"697a6174",
  1209 => x"696f6e20",
  1210 => x"6572726f",
  1211 => x"72210a00",
  1212 => x"434d4435",
  1213 => x"38202564",
  1214 => x"0a202000",
  1215 => x"434d4435",
  1216 => x"385f3220",
  1217 => x"25640a20",
  1218 => x"20000000",
  1219 => x"41637469",
  1220 => x"76617469",
  1221 => x"6e672043",
  1222 => x"530a0000",
  1223 => x"53656e74",
  1224 => x"20726573",
  1225 => x"65742063",
  1226 => x"6f6d6d61",
  1227 => x"6e640a00",
  1228 => x"53442063",
  1229 => x"61726420",
  1230 => x"696e6974",
  1231 => x"69616c69",
  1232 => x"7a617469",
  1233 => x"6f6e2065",
  1234 => x"72726f72",
  1235 => x"210a0000",
  1236 => x"43617264",
  1237 => x"20726573",
  1238 => x"706f6e64",
  1239 => x"65642074",
  1240 => x"6f207265",
  1241 => x"7365740a",
  1242 => x"00000000",
  1243 => x"53444843",
  1244 => x"20636172",
  1245 => x"64206465",
  1246 => x"74656374",
  1247 => x"65640a00",
  1248 => x"53656e64",
  1249 => x"696e6720",
  1250 => x"636d6431",
  1251 => x"360a0000",
  1252 => x"496e6974",
  1253 => x"20646f6e",
  1254 => x"650a0000",
  1255 => x"73645f72",
  1256 => x"6561645f",
  1257 => x"73656374",
  1258 => x"6f722025",
  1259 => x"642c2025",
  1260 => x"640a0000",
  1261 => x"52656164",
  1262 => x"20636f6d",
  1263 => x"6d616e64",
  1264 => x"20666169",
  1265 => x"6c656420",
  1266 => x"61742025",
  1267 => x"64202825",
  1268 => x"64290a00",
  1269 => x"496e6974",
  1270 => x"69616c69",
  1271 => x"7a696e67",
  1272 => x"20534420",
  1273 => x"63617264",
  1274 => x"0a000000",
  1275 => x"48756e74",
  1276 => x"696e6720",
  1277 => x"666f7220",
  1278 => x"70617274",
  1279 => x"6974696f",
  1280 => x"6e0a0000",
  1281 => x"4f53445a",
  1282 => x"50553031",
  1283 => x"53595300",
  1284 => x"43616e27",
  1285 => x"74206c6f",
  1286 => x"61642066",
  1287 => x"69726d77",
  1288 => x"6172650a",
  1289 => x"00000000",
  1290 => x"4661696c",
  1291 => x"65642074",
  1292 => x"6f20696e",
  1293 => x"69746961",
  1294 => x"6c697a65",
  1295 => x"20534420",
  1296 => x"63617264",
  1297 => x"0a000000",
  1298 => x"52656164",
  1299 => x"696e6720",
  1300 => x"4d42520a",
  1301 => x"00000000",
  1302 => x"52656164",
  1303 => x"206f6620",
  1304 => x"4d425220",
  1305 => x"6661696c",
  1306 => x"65640a00",
  1307 => x"4d425220",
  1308 => x"73756363",
  1309 => x"65737366",
  1310 => x"756c6c79",
  1311 => x"20726561",
  1312 => x"640a0000",
  1313 => x"46415431",
  1314 => x"36202020",
  1315 => x"00000000",
  1316 => x"46415433",
  1317 => x"32202020",
  1318 => x"00000000",
  1319 => x"50617274",
  1320 => x"6974696f",
  1321 => x"6e636f75",
  1322 => x"6e742025",
  1323 => x"640a0000",
  1324 => x"4e6f2070",
  1325 => x"61727469",
  1326 => x"74696f6e",
  1327 => x"20736967",
  1328 => x"6e617475",
  1329 => x"72652066",
  1330 => x"6f756e64",
  1331 => x"0a000000",
  1332 => x"52656164",
  1333 => x"696e6720",
  1334 => x"626f6f74",
  1335 => x"20736563",
  1336 => x"746f7220",
  1337 => x"25640a00",
  1338 => x"52656164",
  1339 => x"20626f6f",
  1340 => x"74207365",
  1341 => x"63746f72",
  1342 => x"2066726f",
  1343 => x"6d206669",
  1344 => x"72737420",
  1345 => x"70617274",
  1346 => x"6974696f",
  1347 => x"6e0a0000",
  1348 => x"48756e74",
  1349 => x"696e6720",
  1350 => x"666f7220",
  1351 => x"66696c65",
  1352 => x"73797374",
  1353 => x"656d0a00",
  1354 => x"556e7375",
  1355 => x"70706f72",
  1356 => x"74656420",
  1357 => x"70617274",
  1358 => x"6974696f",
  1359 => x"6e207479",
  1360 => x"7065210d",
  1361 => x"00000000",
  1362 => x"52656164",
  1363 => x"696e6720",
  1364 => x"64697265",
  1365 => x"63746f72",
  1366 => x"79207365",
  1367 => x"63746f72",
  1368 => x"2025640a",
  1369 => x"00000000",
  1370 => x"66696c65",
  1371 => x"20222573",
  1372 => x"2220666f",
  1373 => x"756e640d",
  1374 => x"00000000",
  1375 => x"47657446",
  1376 => x"41544c69",
  1377 => x"6e6b2072",
  1378 => x"65747572",
  1379 => x"6e656420",
  1380 => x"25640a00",
  1381 => x"4f70656e",
  1382 => x"65642066",
  1383 => x"696c652c",
  1384 => x"206c6f61",
  1385 => x"64696e67",
  1386 => x"2e2e2e0a",
  1387 => x"00000000",
  1388 => x"43616e27",
  1389 => x"74206f70",
  1390 => x"656e2025",
  1391 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

